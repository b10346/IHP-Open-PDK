########################################################################
#
# Copyright 2025 IHP PDK Authors
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#    https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
########################################################################

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        0.48 BY 3.78 ;
END  CoreSite

MACRO sg13g2_a21o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21o_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.76 0.405 3.11 0.965 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 1.525 2.545 2 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.525 2.05 2 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6159 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.885 1.225 1.145 ;
        RECT 0.205 2.095 0.56 3.16 ;
        RECT 0.205 0.885 0.445 3.16 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.405 2.585 2.665 4 ;
        RECT 0.81 2.14 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.92 1.145 3.165 1.41 ;
        RECT 2.415 1.145 3.165 1.31 ;
        RECT 2.415 -0.22 2.575 1.31 ;
        RECT 1.455 -0.22 1.715 0.965 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.915 2.21 3.175 3.125 ;
      RECT 1.855 2.21 2.115 3.125 ;
      RECT 1.855 2.21 3.175 2.405 ;
      RECT 1.335 2.17 1.595 3.125 ;
      RECT 1.335 1.54 1.575 3.125 ;
      RECT 1.415 1.145 1.575 3.125 ;
      RECT 0.625 1.54 1.575 1.87 ;
      RECT 1.415 1.145 2.235 1.305 ;
      RECT 2.02 0.825 2.235 1.305 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21o_1

MACRO sg13g2_a21o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21o_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.2 1.56 3.545 2 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.725 1.56 3.02 2 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 1.56 2.535 2 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 2.27 1.08 3.16 ;
        RECT 0.785 0.72 1.045 3.16 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.88 2.55 3.14 4 ;
        RECT 1.295 2.27 1.555 4 ;
        RECT 0.275 2.27 0.535 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.39 -0.22 3.65 1.32 ;
        RECT 1.935 -0.22 2.195 0.99 ;
        RECT 1.295 -0.22 1.555 1.32 ;
        RECT 0.275 -0.22 0.535 1.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 3.39 2.2 3.65 3.16 ;
      RECT 2.33 2.2 2.59 3.16 ;
      RECT 2.33 2.2 3.65 2.36 ;
      RECT 1.81 2.17 2.07 3.16 ;
      RECT 1.81 1.22 2.05 3.16 ;
      RECT 1.235 1.67 2.05 1.93 ;
      RECT 1.81 1.22 2.755 1.38 ;
      RECT 2.495 0.72 2.755 1.38 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21o_2

MACRO sg13g2_a21oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21oi_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.855 -0.22 2.115 1.32 ;
        RECT 0.325 -0.22 0.585 0.98 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.345 2.9 1.605 4 ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.62 1.58 1.88 ;
        RECT 1.32 1.345 1.58 1.88 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.77 1.5 2.115 1.88 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.72 1.095 1.32 ;
        RECT 0.325 2.08 0.995 2.29 ;
        RECT 0.835 0.72 0.995 2.29 ;
        RECT 0.325 2.08 0.62 3.16 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 1.345 0.6 1.88 ;
    END
  END B1
  OBS
    LAYER Metal1 ;
      RECT 1.855 2.08 2.115 3.16 ;
      RECT 0.835 2.555 1.095 3.16 ;
      RECT 0.835 2.555 2.115 2.715 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21oi_1

MACRO sg13g2_a21oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21oi_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.315 -0.22 3.575 1.32 ;
        RECT 2.295 -0.22 2.555 0.98 ;
        RECT 0.255 -0.22 0.515 1.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 1.785 2.95 2.045 4 ;
        RECT 0.765 2.95 1.025 4 ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.24 1.625 3.575 2.28 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.988 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.76 1.16 3.045 2.765 ;
        RECT 2.805 0.72 3.045 2.765 ;
        RECT 1.275 1.16 3.045 1.32 ;
        RECT 1.275 0.785 1.535 1.32 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 2.09 2.3 2.315 ;
        RECT 2.04 1.6 2.3 2.315 ;
        RECT 0.255 1.6 0.77 2.315 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 1.56 1.725 1.9 ;
    END
  END A1
  OBS
    LAYER Metal1 ;
      RECT 2.295 2.965 3.575 3.16 ;
      RECT 3.315 2.56 3.575 3.16 ;
      RECT 1.275 2.565 1.535 3.16 ;
      RECT 0.255 2.565 0.515 3.16 ;
      RECT 2.295 2.565 2.555 3.16 ;
      RECT 0.255 2.565 2.555 2.765 ;
      RECT 0.765 0.445 1.025 1.32 ;
      RECT 1.785 0.445 2.045 0.98 ;
      RECT 0.765 0.445 2.045 0.605 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21oi_2

MACRO sg13g2_a221oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a221oi_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.32 2.505 3.58 4 ;
        RECT 2.3 2.9 2.56 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.32 -0.22 3.58 0.98 ;
        RECT 0.77 -0.22 1.03 0.98 ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 1.555 1.36 1.9 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.555 0.61 1.9 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 1.555 2.04 1.9 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 1.71 2.58 1.94 ;
        RECT 2.26 1.44 2.515 1.94 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1356 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 2.165 3.66 2.325 ;
        RECT 3.5 1.16 3.66 2.325 ;
        RECT 2.81 1.16 3.66 1.37 ;
        RECT 2.81 0.72 3.07 1.37 ;
        RECT 1.28 0.72 3.07 0.98 ;
        RECT 0.26 1.16 1.54 1.37 ;
        RECT 1.28 0.72 1.54 1.37 ;
        RECT 0.26 2.165 0.52 3.16 ;
        RECT 0.26 0.72 0.52 1.37 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 1.57 3.32 1.9 ;
        RECT 2.76 1.57 3.32 1.8 ;
    END
  END A2
  OBS
    LAYER Metal1 ;
      RECT 2.81 2.505 3.07 3.16 ;
      RECT 1.28 2.505 1.54 2.765 ;
      RECT 1.28 2.505 3.07 2.715 ;
      RECT 0.77 2.95 2.05 3.16 ;
      RECT 1.79 2.9 2.05 3.16 ;
      RECT 0.77 2.56 1.03 3.16 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a221oi_1

MACRO sg13g2_a22oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a22oi_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 0.84 1.75 1.1 ;
        RECT 1.31 2.3 1.6 2.9 ;
        RECT 1.42 0.84 1.6 2.9 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.785 1.24 2.07 ;
        RECT 0.82 1.785 1.115 2.255 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 1.77 2.08 2.44 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.33 2.72 2.07 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 1.33 2.09 1.56 ;
        RECT 1.93 0.48 2.09 1.56 ;
        RECT 0.62 0.48 2.09 0.64 ;
        RECT 0.62 0.48 0.78 1.49 ;
        RECT 0.17 1.56 0.64 2.07 ;
        RECT 0.42 1.33 0.64 2.07 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.44 2.3 2.7 4 ;
        RECT 0.18 2.3 0.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.44 -0.22 2.7 1.1 ;
        RECT 0.18 -0.22 0.44 1.1 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.8 3.085 2.08 3.28 ;
      RECT 1.82 2.68 2.08 3.28 ;
      RECT 0.8 2.68 1.06 3.28 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a22oi_1

MACRO sg13g2_and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and2_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.105 0.405 0.78 0.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.435 1.17 1.87 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 2.14 2.275 3.16 ;
        RECT 2.04 0.72 2.275 3.16 ;
        RECT 1.775 0.72 2.275 1.32 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.265 2.56 1.525 4 ;
        RECT 0.245 2.56 0.505 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.265 -0.22 1.525 1.155 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.755 2.05 1.015 3.16 ;
      RECT 0.245 2.05 1.56 2.24 ;
      RECT 1.4 1.605 1.56 2.24 ;
      RECT 0.245 1.14 0.505 2.24 ;
      RECT 1.4 1.605 1.74 1.865 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and2_1

MACRO sg13g2_and2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.105 0.405 0.78 0.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.47 1.17 1.87 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 2.22 2.105 3.16 ;
        RECT 1.92 0.72 2.105 3.16 ;
        RECT 1.775 0.72 2.105 1.32 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.285 2.22 2.545 4 ;
        RECT 1.265 2.56 1.525 4 ;
        RECT 0.245 2.56 0.505 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.285 -0.22 2.545 1.32 ;
        RECT 1.265 -0.22 1.525 1.145 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.755 2.05 1.015 3.16 ;
      RECT 0.245 2.05 1.56 2.24 ;
      RECT 1.4 1.57 1.56 2.24 ;
      RECT 0.245 1.14 0.505 2.24 ;
      RECT 1.4 1.57 1.74 1.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and2_2

MACRO sg13g2_and3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and3_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.78 2.235 3.065 3.175 ;
        RECT 2.895 1.125 3.065 3.175 ;
        RECT 2.44 1.125 3.065 1.385 ;
        RECT 2.44 0.77 2.7 1.385 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.475 1.59 1.09 ;
        RECT 0.35 0.475 1.59 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.4 1.56 1.98 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.4 2.06 1.95 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 1.93 2.575 2.53 4 ;
        RECT 0.91 2.57 1.17 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 1.93 -0.22 2.19 1.14 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.42 2.16 1.68 3.175 ;
      RECT 0.4 1.09 0.66 3.175 ;
      RECT 0.4 2.16 2.405 2.32 ;
      RECT 2.245 1.57 2.405 2.32 ;
      RECT 2.245 1.57 2.645 1.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and3_1

MACRO sg13g2_and3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and3_2 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 2.51 3.02 2.69 ;
        RECT 2.74 1.29 3.02 2.69 ;
        RECT 2.44 1.29 3.02 1.55 ;
        RECT 2.435 2.51 2.705 3.175 ;
        RECT 2.44 0.77 2.7 1.55 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.475 1.59 1.09 ;
        RECT 0.35 0.475 1.59 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.125 1.4 1.56 1.95 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.76 1.4 2.06 1.95 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.95 2.915 3.21 4 ;
        RECT 1.93 2.575 2.19 4 ;
        RECT 0.91 2.575 1.17 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.95 -0.22 3.21 1.09 ;
        RECT 1.93 -0.22 2.19 1.14 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.415 2.16 1.675 3.175 ;
      RECT 0.4 1.09 0.66 3.175 ;
      RECT 0.4 2.16 2.43 2.32 ;
      RECT 2.27 1.77 2.43 2.32 ;
      RECT 2.27 1.77 2.53 2.03 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and3_2

MACRO sg13g2_and4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and4_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.725 1.455 1.08 1.985 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 1.455 1.56 1.985 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 1.455 2.045 1.985 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 1.45 2.665 2 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8928 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 2.07 3.685 3.18 ;
        RECT 3.525 0.61 3.685 3.18 ;
        RECT 3.205 0.61 3.685 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.54 2.56 2.8 4 ;
        RECT 1.445 2.56 1.705 4 ;
        RECT 0.425 2.56 0.685 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.55 -0.22 2.815 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.935 2.22 1.195 3.125 ;
      RECT 1.985 2.22 2.245 3.12 ;
      RECT 0.355 2.22 3.01 2.38 ;
      RECT 2.85 1.54 3.01 2.38 ;
      RECT 0.355 0.61 0.525 2.38 ;
      RECT 2.85 1.54 3.205 1.87 ;
      RECT 0.355 0.61 0.685 1.21 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and4_1

MACRO sg13g2_and4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and4_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.765 1.35 1.08 2.01 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.285 1.35 1.565 2.01 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 1.35 2.06 2.01 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.28 1.46 2.615 2.01 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 2.21 3.685 3.16 ;
        RECT 3.525 0.64 3.685 3.16 ;
        RECT 3.205 0.64 3.685 1.26 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.865 2.21 4.125 4 ;
        RECT 2.54 2.56 2.8 4 ;
        RECT 1.445 2.56 1.705 4 ;
        RECT 0.425 2.56 0.685 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.865 -0.22 4.125 1.21 ;
        RECT 2.55 -0.22 2.815 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.985 2.22 2.245 3.16 ;
      RECT 0.935 2.22 1.195 3.16 ;
      RECT 0.265 2.22 3.01 2.38 ;
      RECT 2.85 1.54 3.01 2.38 ;
      RECT 0.265 0.645 0.435 2.38 ;
      RECT 2.85 1.54 3.205 1.87 ;
      RECT 0.265 0.645 0.685 1.17 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and4_2

MACRO sg13g2_antennanp
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_antennanp 0 0 ;
  SIZE 1.44 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.44 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.44 0.22 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0154 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.57 1.05 1.16 ;
        RECT 0.38 2.08 0.98 2.68 ;
        RECT 0.38 1.13 0.63 2.68 ;
    END
  END A
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_antennanp

MACRO sg13g2_buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1.93 0.68 2.26 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 2.02 1.6 3.18 ;
        RECT 1.41 0.55 1.6 3.18 ;
        RECT 1.31 0.55 1.6 1.29 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.77 2.89 1.03 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.765 -0.22 1.015 1.07 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.24 2.44 0.51 3.18 ;
      RECT 0.24 2.44 1.07 2.62 ;
      RECT 0.9 1.29 1.07 2.62 ;
      RECT 0.9 1.5 1.225 1.83 ;
      RECT 0.215 1.29 1.07 1.465 ;
      RECT 0.215 1 0.515 1.465 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_1

MACRO sg13g2_buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_16 0 0 ;
  SIZE 12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.6544 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.91 2.2 8.17 3.16 ;
        RECT 5.87 1.05 8.17 1.22 ;
        RECT 7.91 0.61 8.17 1.22 ;
        RECT 2.81 2.2 8.17 2.36 ;
        RECT 6.89 2.2 7.15 3.16 ;
        RECT 6.89 0.61 7.15 1.22 ;
        RECT 5.87 0.61 6.13 3.16 ;
        RECT 4.85 0.61 5.11 3.16 ;
        RECT 3.83 0.61 4.09 3.16 ;
        RECT 2.81 0.61 3.07 3.16 ;
        RECT 1.79 1.52 3.07 1.85 ;
        RECT 1.79 0.61 2.05 3.16 ;
        RECT 0.77 2.2 2.05 2.36 ;
        RECT 0.77 0.61 1.03 3.16 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4508 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.26 1.52 11.44 1.85 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12 4 ;
        RECT 11.48 2.215 11.74 4 ;
        RECT 10.46 2.545 10.72 4 ;
        RECT 9.44 2.54 9.7 4 ;
        RECT 8.42 2.54 8.68 4 ;
        RECT 7.4 2.54 7.66 4 ;
        RECT 6.38 2.54 6.64 4 ;
        RECT 5.36 2.54 5.62 4 ;
        RECT 4.34 2.54 4.6 4 ;
        RECT 3.32 2.54 3.58 4 ;
        RECT 2.3 2.22 2.56 4 ;
        RECT 1.28 2.54 1.54 4 ;
        RECT 0.26 2.22 0.52 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12 0.22 ;
        RECT 11.48 -0.22 11.74 1.21 ;
        RECT 10.46 -0.22 10.72 0.87 ;
        RECT 9.44 -0.22 9.7 0.87 ;
        RECT 8.42 -0.22 8.685 0.87 ;
        RECT 7.4 -0.22 7.66 0.87 ;
        RECT 6.38 -0.22 6.64 0.87 ;
        RECT 5.36 -0.22 5.62 1.195 ;
        RECT 4.34 -0.22 4.6 1.195 ;
        RECT 3.32 -0.22 3.58 1.195 ;
        RECT 2.3 -0.22 2.56 1.21 ;
        RECT 1.28 -0.22 1.54 1.21 ;
        RECT 0.26 -0.22 0.52 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 10.97 2.2 11.23 3.16 ;
      RECT 9.95 2.2 10.21 3.16 ;
      RECT 8.93 2.2 9.19 3.16 ;
      RECT 8.385 2.2 11.23 2.36 ;
      RECT 8.385 1.05 8.595 2.36 ;
      RECT 6.395 1.52 8.595 1.85 ;
      RECT 8.385 1.05 11.23 1.22 ;
      RECT 10.97 0.61 11.23 1.22 ;
      RECT 9.95 0.61 10.21 1.22 ;
      RECT 8.93 0.61 9.19 1.22 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_16

MACRO sg13g2_buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_2 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.49 2.14 1.87 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 0.61 1.235 2.34 ;
        RECT 0.67 1.52 1.235 1.85 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.485 2.895 1.745 4 ;
        RECT 0.15 2.56 0.41 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.485 -0.22 1.745 0.965 ;
        RECT 0.465 -0.22 0.725 1.31 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.97 2.18 2.26 3.1 ;
      RECT 0.605 2.55 2.26 2.71 ;
      RECT 1.415 1.145 1.575 2.71 ;
      RECT 0.605 2.215 0.765 2.71 ;
      RECT 0.225 2.215 0.765 2.375 ;
      RECT 0.225 1.555 0.485 2.375 ;
      RECT 1.415 1.145 2.255 1.31 ;
      RECT 1.995 0.72 2.255 1.31 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_2

MACRO sg13g2_buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_4 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.995 2.025 3.13 ;
        RECT 0.745 1.065 2.025 1.225 ;
        RECT 1.765 0.645 2.025 1.225 ;
        RECT 0.745 1.995 2.025 2.165 ;
        RECT 0.745 0.605 1.005 3.13 ;
        RECT 0.32 1.525 1.005 1.84 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 1.475 3.15 1.885 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.295 2.64 3.555 4 ;
        RECT 2.275 2.08 2.535 4 ;
        RECT 1.255 2.49 1.515 4 ;
        RECT 0.235 2.115 0.495 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.375 0.61 2.975 0.87 ;
        RECT 2.545 -0.22 2.805 0.87 ;
        RECT 1.255 -0.22 1.515 0.87 ;
        RECT 0.235 -0.22 0.495 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.785 2.15 3.045 2.77 ;
      RECT 2.785 2.15 3.59 2.42 ;
      RECT 3.4 0.64 3.59 2.42 ;
      RECT 1.68 1.54 2.43 1.8 ;
      RECT 2.265 1.05 2.43 1.8 ;
      RECT 2.265 1.05 3.59 1.21 ;
      RECT 3.245 0.64 3.59 1.21 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_4

MACRO sg13g2_buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_8 0 0 ;
  SIZE 6.24 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.7254 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 1.5 1.51 1.865 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 1.55 5.95 1.815 ;
        RECT 5.26 0.61 5.52 3.16 ;
        RECT 2.2 2.22 5.52 2.38 ;
        RECT 2.2 1.05 5.52 1.21 ;
        RECT 4.24 2.22 4.5 3.16 ;
        RECT 4.24 0.61 4.5 1.21 ;
        RECT 3.22 2.22 3.48 3.16 ;
        RECT 3.22 0.61 3.48 1.21 ;
        RECT 2.2 2.22 2.46 3.16 ;
        RECT 2.2 0.61 2.46 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 6.24 4 ;
        RECT 5.77 2.22 6.03 4 ;
        RECT 4.75 2.56 5.01 4 ;
        RECT 3.73 2.56 3.99 4 ;
        RECT 2.71 2.56 2.97 4 ;
        RECT 1.69 2.56 1.95 4 ;
        RECT 0.67 2.56 0.93 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 6.24 0.22 ;
        RECT 5.77 -0.22 6.03 1.21 ;
        RECT 4.75 -0.22 5.01 0.87 ;
        RECT 3.73 -0.22 3.99 0.87 ;
        RECT 2.71 -0.22 2.97 0.87 ;
        RECT 1.69 -0.22 1.95 0.87 ;
        RECT 0.67 -0.22 0.93 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.18 2.22 1.44 3.16 ;
      RECT 0.16 2.22 0.42 3.16 ;
      RECT 0.16 2.22 1.94 2.38 ;
      RECT 1.77 1.05 1.94 2.38 ;
      RECT 1.77 1.555 4.975 1.815 ;
      RECT 0.16 1.05 1.94 1.21 ;
      RECT 1.18 0.61 1.44 1.21 ;
      RECT 0.16 0.61 0.42 1.21 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_8

MACRO sg13g2_decap_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_decap_4 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.065 2.22 1.79 4 ;
        RECT 1.065 1.47 1.405 4 ;
        RECT 0.13 2.22 0.4 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.51 -0.22 1.79 0.935 ;
        RECT 0.53 -0.22 0.855 1.805 ;
        RECT 0.13 -0.22 0.855 0.935 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_decap_4

MACRO sg13g2_decap_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_decap_8 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.945 2.21 3.205 4 ;
        RECT 1.22 1.475 2.155 4 ;
        RECT 0.185 2.205 0.445 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.585 -0.22 3.195 0.99 ;
        RECT 2.585 -0.22 2.835 1.81 ;
        RECT 1.53 -0.22 1.835 1.03 ;
        RECT 0.52 -0.22 0.81 1.81 ;
        RECT 0.175 -0.22 0.81 0.99 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_decap_8

MACRO sg13g2_dfrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbp_1 0 0 ;
  SIZE 13.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8998 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.746642 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.145 1.51 2.75 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 13.92 0.22 ;
        RECT 12.635 -0.22 12.895 1.19 ;
        RECT 10.91 -0.22 11.15 0.85 ;
        RECT 9.56 -0.22 9.82 0.85 ;
        RECT 2.235 -0.22 2.495 0.915 ;
        RECT 1.14 -0.22 1.41 0.85 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 13.92 4 ;
        RECT 12.63 2.1 12.9 4 ;
        RECT 10.89 2.46 11.15 4 ;
        RECT 2.945 2.86 3.115 4 ;
        RECT 0.215 2.24 0.475 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1.07 0.6 1.89 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.145 2.095 13.56 3.155 ;
        RECT 13.35 0.59 13.56 3.155 ;
        RECT 13.125 0.59 13.56 1.19 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7161 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.34 0.99 11.725 1.52 ;
        RECT 11.4 0.59 11.66 3.155 ;
    END
  END Q_N
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.45 1.52 6.99 1.84 ;
    END
  END CLK
  OBS
    LAYER Metal1 ;
      RECT 12.125 0.59 12.385 3.155 ;
      RECT 12.87 1.445 13.17 1.745 ;
      RECT 12.125 1.485 13.17 1.71 ;
      RECT 10.07 2.035 10.33 2.495 ;
      RECT 9.22 2.035 11 2.195 ;
      RECT 10.84 1.03 11 2.195 ;
      RECT 9.22 1.69 9.48 2.195 ;
      RECT 10.57 1.03 11 1.19 ;
      RECT 10.57 0.625 10.73 1.19 ;
      RECT 10.38 0.625 10.73 0.885 ;
      RECT 8.475 2.225 8.95 2.485 ;
      RECT 8.79 1.145 8.95 2.485 ;
      RECT 10.165 1.35 10.47 1.625 ;
      RECT 8.79 1.35 10.47 1.51 ;
      RECT 8.79 1.145 8.97 1.51 ;
      RECT 7.96 1.145 8.97 1.315 ;
      RECT 9.91 3.025 10.16 3.285 ;
      RECT 4.855 3.025 5.115 3.285 ;
      RECT 4.855 3.075 10.16 3.235 ;
      RECT 7.51 0.805 7.725 1.31 ;
      RECT 7.51 0.805 9.31 0.965 ;
      RECT 9.05 0.59 9.31 0.965 ;
      RECT 1.2 2.5 1.94 2.76 ;
      RECT 1.2 1.15 1.36 2.76 ;
      RECT 7.745 1.555 7.935 2.425 ;
      RECT 2.95 1.705 3.21 1.965 ;
      RECT 7.17 1.555 7.935 1.725 ;
      RECT 2.95 1.15 3.11 1.965 ;
      RECT 7.17 0.44 7.33 1.725 ;
      RECT 1.2 1.15 3.11 1.31 ;
      RECT 2.705 0.44 2.875 1.31 ;
      RECT 1.72 0.815 1.98 1.31 ;
      RECT 8.54 0.44 8.8 0.625 ;
      RECT 2.705 0.44 8.8 0.605 ;
      RECT 5.55 2.63 8.275 2.8 ;
      RECT 8.115 1.525 8.275 2.8 ;
      RECT 5.55 2.07 5.81 2.8 ;
      RECT 4.855 2.16 5.81 2.42 ;
      RECT 5.145 2.07 5.81 2.42 ;
      RECT 5.145 0.92 5.42 2.42 ;
      RECT 8.115 1.525 8.6 1.785 ;
      RECT 5.145 0.92 5.815 1.18 ;
      RECT 6.02 2.07 7.525 2.33 ;
      RECT 6.02 0.98 6.18 2.33 ;
      RECT 5.725 1.575 6.18 1.835 ;
      RECT 6.755 0.92 6.99 1.18 ;
      RECT 6.02 0.98 6.99 1.14 ;
      RECT 4.66 1.44 4.905 1.7 ;
      RECT 4.725 0.785 4.905 1.7 ;
      RECT 3.12 0.785 4.905 0.96 ;
      RECT 3.365 3.08 4.505 3.24 ;
      RECT 4.32 2.655 4.505 3.24 ;
      RECT 0.785 3.08 2.765 3.24 ;
      RECT 2.605 2.52 2.765 3.24 ;
      RECT 3.365 2.52 3.535 3.24 ;
      RECT 0.785 0.59 0.95 3.24 ;
      RECT 4.32 2.655 4.665 2.915 ;
      RECT 2.605 2.52 3.535 2.68 ;
      RECT 4.32 1.16 4.48 3.24 ;
      RECT 0.72 2.24 0.98 2.5 ;
      RECT 3.385 1.16 3.645 1.64 ;
      RECT 3.385 1.16 4.48 1.32 ;
      RECT 0.21 0.59 0.95 0.85 ;
      RECT 2.245 2.145 2.425 2.9 ;
      RECT 3.895 1.5 4.115 2.805 ;
      RECT 2.245 2.145 4.115 2.315 ;
      RECT 1.585 2.145 4.115 2.305 ;
      RECT 1.585 1.705 1.845 2.305 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbp_1

MACRO sg13g2_dfrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbp_2 0 0 ;
  SIZE 14.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 1.51 2.75 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 14.4 0.22 ;
        RECT 13.935 -0.22 14.21 0.84 ;
        RECT 12.93 -0.22 13.19 1.21 ;
        RECT 11.91 -0.22 12.17 0.85 ;
        RECT 10.91 -0.22 11.15 0.85 ;
        RECT 9.56 -0.22 9.82 0.885 ;
        RECT 2.235 -0.22 2.495 0.915 ;
        RECT 1.14 -0.22 1.4 0.885 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 14.4 4 ;
        RECT 13.58 2.085 13.84 4 ;
        RECT 12.555 2.085 12.815 4 ;
        RECT 11.47 1.98 11.73 4 ;
        RECT 10.45 2.46 10.71 4 ;
        RECT 2.945 2.86 3.115 4 ;
        RECT 0.215 2.215 0.47 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1.375 0.61 1.855 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7124 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.44 1.045 14.21 1.49 ;
        RECT 13.19 1.515 13.7 1.775 ;
        RECT 13.44 0.595 13.7 1.775 ;
        RECT 13.065 2.085 13.36 3.175 ;
        RECT 13.19 1.515 13.36 3.175 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.96 1.52 11.72 1.74 ;
        RECT 11.34 0.99 11.72 1.74 ;
        RECT 11.395 0.59 11.66 1.74 ;
        RECT 10.96 1.52 11.22 3.06 ;
    END
  END Q_N
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.365 1.335 6.99 1.935 ;
    END
  END CLK
  OBS
    LAYER Metal1 ;
      RECT 11.98 1.98 12.36 2.92 ;
      RECT 12.19 1.535 12.36 2.92 ;
      RECT 12.19 1.535 12.985 1.795 ;
      RECT 12.4 0.59 12.685 1.795 ;
      RECT 9.91 2.1 10.17 2.495 ;
      RECT 9.13 2.1 10.73 2.26 ;
      RECT 10.57 0.625 10.73 2.26 ;
      RECT 9.13 1.655 9.385 2.26 ;
      RECT 10.38 0.625 10.73 0.885 ;
      RECT 8.455 2.125 8.66 2.5 ;
      RECT 8.455 2.125 8.95 2.295 ;
      RECT 8.79 1.145 8.95 2.295 ;
      RECT 10.165 1.275 10.39 1.665 ;
      RECT 8.79 1.275 10.39 1.465 ;
      RECT 7.96 1.145 8.97 1.315 ;
      RECT 9.91 3.025 10.18 3.285 ;
      RECT 4.855 3.025 5.115 3.285 ;
      RECT 4.855 3.075 10.18 3.235 ;
      RECT 7.51 0.805 7.68 1.31 ;
      RECT 7.51 0.805 9.31 0.965 ;
      RECT 9.05 0.625 9.31 0.965 ;
      RECT 1.2 2.64 1.94 2.9 ;
      RECT 1.2 1.17 1.36 2.9 ;
      RECT 7.745 1.555 7.935 2.45 ;
      RECT 2.935 1.755 3.215 1.965 ;
      RECT 2.935 1.17 3.095 1.965 ;
      RECT 7.17 1.555 7.935 1.725 ;
      RECT 7.17 0.44 7.33 1.725 ;
      RECT 1.2 1.17 3.095 1.33 ;
      RECT 2.705 0.44 2.875 1.33 ;
      RECT 1.72 0.815 1.98 1.33 ;
      RECT 8.54 0.44 8.8 0.625 ;
      RECT 2.705 0.44 8.8 0.605 ;
      RECT 5.425 2.63 8.275 2.79 ;
      RECT 8.115 1.51 8.275 2.79 ;
      RECT 5.425 2.06 5.785 2.79 ;
      RECT 5.02 2.15 5.785 2.41 ;
      RECT 5.155 2.06 5.785 2.41 ;
      RECT 5.155 1.135 5.415 2.41 ;
      RECT 8.115 1.51 8.6 1.77 ;
      RECT 5.965 2.145 7.525 2.37 ;
      RECT 7.265 2.075 7.525 2.37 ;
      RECT 5.965 0.855 6.125 2.37 ;
      RECT 5.65 1.54 6.125 1.87 ;
      RECT 6.755 0.81 6.99 1.07 ;
      RECT 5.965 0.855 6.99 1.025 ;
      RECT 4.63 1.44 4.895 1.7 ;
      RECT 4.685 1.3 4.895 1.7 ;
      RECT 4.685 0.785 4.865 1.7 ;
      RECT 3.165 0.785 4.865 0.96 ;
      RECT 0.79 3.08 2.765 3.24 ;
      RECT 2.605 2.52 2.765 3.24 ;
      RECT 3.455 2.985 4.625 3.145 ;
      RECT 4.29 2.685 4.625 3.145 ;
      RECT 0.79 2.24 0.98 3.24 ;
      RECT 3.455 2.52 3.615 3.145 ;
      RECT 4.29 1.17 4.45 3.145 ;
      RECT 2.605 2.52 3.615 2.68 ;
      RECT 0.72 2.24 0.98 2.52 ;
      RECT 0.79 0.645 0.95 3.24 ;
      RECT 3.385 1.225 3.645 1.64 ;
      RECT 3.465 1.17 4.45 1.33 ;
      RECT 0.21 0.645 0.95 0.84 ;
      RECT 2.245 2.145 2.425 2.9 ;
      RECT 3.89 1.51 4.075 2.805 ;
      RECT 2.245 2.145 4.075 2.315 ;
      RECT 1.585 2.145 4.075 2.305 ;
      RECT 1.585 1.705 1.845 2.305 ;
      RECT 3.89 1.51 4.11 1.81 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbp_2

MACRO sg13g2_dfrbpq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbpq_1 0 0 ;
  SIZE 12.96 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8998 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.746642 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.145 1.51 2.75 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12.96 0.22 ;
        RECT 11.785 -0.22 12.045 1.19 ;
        RECT 9.56 -0.22 9.82 0.85 ;
        RECT 2.235 -0.22 2.495 0.915 ;
        RECT 1.14 -0.22 1.41 0.85 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12.96 4 ;
        RECT 11.785 2.1 12.045 4 ;
        RECT 10.61 2.225 10.875 4 ;
        RECT 2.945 2.86 3.115 4 ;
        RECT 0.215 2.24 0.475 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1.07 0.6 1.89 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.295 2.095 12.71 3.155 ;
        RECT 12.5 0.59 12.71 3.155 ;
        RECT 12.275 0.59 12.71 1.19 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.45 1.52 6.99 1.84 ;
    END
  END CLK
  OBS
    LAYER Metal1 ;
      RECT 11.275 0.59 11.535 3.155 ;
      RECT 12.02 1.445 12.32 1.745 ;
      RECT 11.275 1.485 12.32 1.71 ;
      RECT 10.07 1.86 10.33 2.495 ;
      RECT 9.22 1.86 10.835 2.02 ;
      RECT 10.675 1.03 10.835 2.02 ;
      RECT 9.22 1.69 9.48 2.02 ;
      RECT 10.57 0.625 10.73 1.19 ;
      RECT 10.38 0.625 10.73 0.885 ;
      RECT 8.475 2.225 8.95 2.485 ;
      RECT 8.79 1.145 8.95 2.485 ;
      RECT 10.165 1.35 10.47 1.625 ;
      RECT 8.79 1.35 10.47 1.51 ;
      RECT 8.79 1.145 8.97 1.51 ;
      RECT 7.96 1.145 8.97 1.315 ;
      RECT 9.91 3.025 10.16 3.285 ;
      RECT 4.855 3.025 5.115 3.285 ;
      RECT 4.855 3.075 10.16 3.235 ;
      RECT 7.51 0.805 7.725 1.31 ;
      RECT 7.51 0.805 9.31 0.965 ;
      RECT 9.05 0.59 9.31 0.965 ;
      RECT 1.2 2.5 1.94 2.76 ;
      RECT 1.2 1.15 1.36 2.76 ;
      RECT 7.745 1.555 7.935 2.425 ;
      RECT 2.95 1.705 3.21 1.965 ;
      RECT 7.17 1.555 7.935 1.725 ;
      RECT 2.95 1.15 3.11 1.965 ;
      RECT 7.17 0.44 7.33 1.725 ;
      RECT 1.2 1.15 3.11 1.31 ;
      RECT 2.705 0.44 2.875 1.31 ;
      RECT 1.72 0.815 1.98 1.31 ;
      RECT 8.54 0.44 8.8 0.625 ;
      RECT 2.705 0.44 8.8 0.605 ;
      RECT 5.55 2.63 8.275 2.8 ;
      RECT 8.115 1.525 8.275 2.8 ;
      RECT 5.55 2.07 5.81 2.8 ;
      RECT 4.855 2.16 5.81 2.42 ;
      RECT 5.145 2.07 5.81 2.42 ;
      RECT 5.145 0.92 5.42 2.42 ;
      RECT 8.115 1.525 8.6 1.785 ;
      RECT 5.145 0.92 5.815 1.18 ;
      RECT 6.02 2.07 7.525 2.33 ;
      RECT 6.02 0.98 6.18 2.33 ;
      RECT 5.725 1.575 6.18 1.835 ;
      RECT 6.755 0.92 6.99 1.18 ;
      RECT 6.02 0.98 6.99 1.14 ;
      RECT 4.66 1.44 4.905 1.7 ;
      RECT 4.725 0.785 4.905 1.7 ;
      RECT 3.12 0.785 4.905 0.96 ;
      RECT 3.365 3.08 4.505 3.24 ;
      RECT 4.32 2.655 4.505 3.24 ;
      RECT 0.785 3.08 2.765 3.24 ;
      RECT 2.605 2.52 2.765 3.24 ;
      RECT 3.365 2.52 3.535 3.24 ;
      RECT 0.785 0.59 0.95 3.24 ;
      RECT 4.32 2.655 4.665 2.915 ;
      RECT 2.605 2.52 3.535 2.68 ;
      RECT 4.32 1.16 4.48 3.24 ;
      RECT 0.72 2.24 0.98 2.5 ;
      RECT 3.385 1.16 3.645 1.64 ;
      RECT 3.385 1.16 4.48 1.32 ;
      RECT 0.21 0.59 0.95 0.85 ;
      RECT 2.245 2.145 2.425 2.9 ;
      RECT 3.895 1.5 4.115 2.805 ;
      RECT 2.245 2.145 4.115 2.315 ;
      RECT 1.585 2.145 4.115 2.305 ;
      RECT 1.585 1.705 1.845 2.305 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbpq_1

MACRO sg13g2_dfrbpq_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbpq_2 0 0 ;
  SIZE 13.44 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 1.51 2.75 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 13.44 0.22 ;
        RECT 12.96 -0.22 13.215 1.2 ;
        RECT 11.935 -0.22 12.2 1.2 ;
        RECT 10.925 -0.22 11.16 1.19 ;
        RECT 9.56 -0.22 9.82 0.885 ;
        RECT 2.235 -0.22 2.495 0.915 ;
        RECT 1.14 -0.22 1.4 0.885 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 13.44 4 ;
        RECT 12.955 2.22 13.215 4 ;
        RECT 11.93 2.19 12.19 4 ;
        RECT 10.45 2.46 10.71 4 ;
        RECT 2.945 2.86 3.115 4 ;
        RECT 0.215 2.215 0.47 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1.375 0.61 1.855 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7161 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.44 1.505 13.15 1.845 ;
        RECT 12.44 0.595 12.7 3.16 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.365 1.335 6.99 1.935 ;
    END
  END CLK
  OBS
    LAYER Metal1 ;
      RECT 10.99 1.555 11.25 3.105 ;
      RECT 10.99 1.555 11.92 1.795 ;
      RECT 11.41 1.54 11.92 1.795 ;
      RECT 11.41 0.59 11.67 1.795 ;
      RECT 9.91 2.1 10.17 2.495 ;
      RECT 9.13 2.1 10.73 2.26 ;
      RECT 10.57 0.625 10.73 2.26 ;
      RECT 9.13 1.655 9.385 2.26 ;
      RECT 10.38 0.625 10.73 0.885 ;
      RECT 8.455 2.125 8.66 2.5 ;
      RECT 8.455 2.125 8.95 2.295 ;
      RECT 8.79 1.145 8.95 2.295 ;
      RECT 10.165 1.275 10.39 1.665 ;
      RECT 8.79 1.275 10.39 1.465 ;
      RECT 7.96 1.145 8.97 1.315 ;
      RECT 9.91 3.025 10.18 3.285 ;
      RECT 4.855 3.025 5.115 3.285 ;
      RECT 4.855 3.075 10.18 3.235 ;
      RECT 7.51 0.805 7.68 1.31 ;
      RECT 7.51 0.805 9.31 0.965 ;
      RECT 9.05 0.625 9.31 0.965 ;
      RECT 1.2 2.64 1.94 2.9 ;
      RECT 1.2 1.17 1.36 2.9 ;
      RECT 7.745 1.555 7.935 2.45 ;
      RECT 2.935 1.755 3.215 1.965 ;
      RECT 2.935 1.17 3.095 1.965 ;
      RECT 7.17 1.555 7.935 1.725 ;
      RECT 7.17 0.44 7.33 1.725 ;
      RECT 1.2 1.17 3.095 1.33 ;
      RECT 2.705 0.44 2.875 1.33 ;
      RECT 1.72 0.815 1.98 1.33 ;
      RECT 8.54 0.44 8.8 0.625 ;
      RECT 2.705 0.44 8.8 0.605 ;
      RECT 5.425 2.63 8.275 2.79 ;
      RECT 8.115 1.51 8.275 2.79 ;
      RECT 5.425 2.06 5.785 2.79 ;
      RECT 5.02 2.15 5.785 2.41 ;
      RECT 5.155 2.06 5.785 2.41 ;
      RECT 5.155 1.135 5.415 2.41 ;
      RECT 8.115 1.51 8.6 1.77 ;
      RECT 5.965 2.145 7.525 2.37 ;
      RECT 7.265 2.075 7.525 2.37 ;
      RECT 5.965 0.855 6.125 2.37 ;
      RECT 5.65 1.54 6.125 1.87 ;
      RECT 6.755 0.81 6.99 1.07 ;
      RECT 5.965 0.855 6.99 1.025 ;
      RECT 4.63 1.44 4.895 1.7 ;
      RECT 4.685 1.3 4.895 1.7 ;
      RECT 4.685 0.785 4.865 1.7 ;
      RECT 3.165 0.785 4.865 0.96 ;
      RECT 0.79 3.08 2.765 3.24 ;
      RECT 2.605 2.52 2.765 3.24 ;
      RECT 3.455 2.985 4.625 3.145 ;
      RECT 4.29 2.685 4.625 3.145 ;
      RECT 0.79 2.24 0.98 3.24 ;
      RECT 3.455 2.52 3.615 3.145 ;
      RECT 4.29 1.17 4.45 3.145 ;
      RECT 2.605 2.52 3.615 2.68 ;
      RECT 0.72 2.24 0.98 2.52 ;
      RECT 0.79 0.645 0.95 3.24 ;
      RECT 3.385 1.225 3.645 1.64 ;
      RECT 3.465 1.17 4.45 1.33 ;
      RECT 0.21 0.645 0.95 0.84 ;
      RECT 2.245 2.145 2.425 2.9 ;
      RECT 3.89 1.51 4.075 2.805 ;
      RECT 2.245 2.145 4.075 2.315 ;
      RECT 1.585 2.145 4.075 2.305 ;
      RECT 1.585 1.705 1.845 2.305 ;
      RECT 3.89 1.51 4.11 1.81 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbpq_2

MACRO sg13g2_dlhq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhq_1 0 0 ;
  SIZE 8.16 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.315 1.4 0.785 2.07 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.575 1.57 6.905 2 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.45 2.075 7.785 3.155 ;
        RECT 7.625 0.63 7.785 3.155 ;
        RECT 7.435 0.63 7.785 1.355 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.16 4 ;
        RECT 6.965 2.23 7.225 4 ;
        RECT 5.03 3.115 5.305 4 ;
        RECT 1.85 3.19 2.11 4 ;
        RECT 0.275 2.4 0.535 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.16 0.22 ;
        RECT 6.88 -0.22 7.14 0.515 ;
        RECT 5.27 -0.22 5.55 0.445 ;
        RECT 1.925 -0.22 2.185 1.27 ;
        RECT 0.335 -0.22 0.595 1.03 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 4.5 1.93 5.005 2.195 ;
      RECT 4.77 0.475 5.005 2.195 ;
      RECT 7.085 1.54 7.445 1.87 ;
      RECT 7.085 0.7 7.255 1.87 ;
      RECT 6.29 0.7 7.255 0.88 ;
      RECT 4.77 0.625 6.5 0.785 ;
      RECT 2.39 0.475 2.665 0.78 ;
      RECT 2.39 0.475 5.005 0.635 ;
      RECT 3.78 2.725 6.715 2.885 ;
      RECT 6.035 2.205 6.715 2.885 ;
      RECT 3.78 1.93 3.95 2.885 ;
      RECT 6.035 1.57 6.395 2.885 ;
      RECT 6.235 1.115 6.395 2.885 ;
      RECT 3.39 1.93 3.95 2.095 ;
      RECT 3.045 1.655 3.545 1.975 ;
      RECT 6.235 1.115 6.6 1.39 ;
      RECT 4.13 2.385 5.815 2.545 ;
      RECT 5.565 1.005 5.815 2.545 ;
      RECT 4.13 1.515 4.29 2.545 ;
      RECT 3.735 1.515 4.29 1.75 ;
      RECT 5.565 1.005 6.055 1.265 ;
      RECT 3.05 2.275 3.6 2.435 ;
      RECT 2.705 2.155 3.205 2.315 ;
      RECT 2.705 1.315 2.865 2.315 ;
      RECT 2.705 1.315 3.545 1.475 ;
      RECT 4.255 0.995 4.585 1.325 ;
      RECT 3.225 1.155 4.585 1.325 ;
      RECT 3.33 3.065 4.175 3.235 ;
      RECT 3.33 2.615 3.5 3.235 ;
      RECT 2.71 2.615 3.5 2.785 ;
      RECT 2.27 2.495 2.865 2.66 ;
      RECT 2.27 2.225 2.52 2.66 ;
      RECT 1.535 1.575 2.525 1.745 ;
      RECT 2.365 0.965 2.525 1.745 ;
      RECT 1.535 0.725 1.695 1.745 ;
      RECT 2.365 0.965 3.02 1.13 ;
      RECT 1.415 0.725 1.695 1.035 ;
      RECT 2.85 0.815 4.02 0.975 ;
      RECT 2.355 3.025 3.04 3.205 ;
      RECT 1.335 2.215 1.57 3.165 ;
      RECT 2.355 2.84 2.525 3.205 ;
      RECT 1.335 2.84 2.525 3 ;
      RECT 0.785 2.405 1.135 3.135 ;
      RECT 0.965 1.32 1.135 3.135 ;
      RECT 0.965 1.32 1.355 1.99 ;
      RECT 0.965 0.79 1.125 3.135 ;
      RECT 0.825 0.79 1.125 1.095 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhq_1

MACRO sg13g2_dlhr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhr_1 0 0 ;
  SIZE 8.64 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.765 1.45 1.11 1.91 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.29 1.45 1.59 1.91 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.63 1.325 6.05 1.875 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.53 2.395 6.945 3.175 ;
        RECT 6.785 1.01 6.945 3.175 ;
        RECT 6.435 1.01 6.945 1.24 ;
        RECT 6.435 0.51 6.72 1.24 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.64 4 ;
        RECT 7.635 2.31 7.82 4 ;
        RECT 6.095 2.46 6.285 4 ;
        RECT 4.7 2.835 5.3 4 ;
        RECT 2.65 2.935 2.93 4 ;
        RECT 0.97 2.935 1.23 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.64 0.22 ;
        RECT 7.55 -0.22 7.81 1.12 ;
        RECT 5.905 -0.22 6.235 1.14 ;
        RECT 4.545 -0.22 4.83 1.115 ;
        RECT 2.645 -0.22 2.905 0.54 ;
        RECT 0.91 -0.22 1.24 1.25 ;
    END
  END VSS
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8 1.97 8.39 3.09 ;
        RECT 8.215 0.47 8.39 3.09 ;
        RECT 8.02 0.47 8.39 1.085 ;
    END
  END Q_N
  OBS
    LAYER Metal1 ;
      RECT 7.125 1.475 7.315 3.09 ;
      RECT 7.125 1.475 8 1.76 ;
      RECT 7.125 0.49 7.305 3.09 ;
      RECT 7 0.49 7.305 0.775 ;
      RECT 5.575 2.055 5.78 3.09 ;
      RECT 4.51 2.12 5.78 2.45 ;
      RECT 6.29 1.48 6.605 2.215 ;
      RECT 5.29 2.055 6.605 2.215 ;
      RECT 5.29 0.51 5.45 2.45 ;
      RECT 5.085 0.51 5.45 1.23 ;
      RECT 3.495 2.535 3.8 2.855 ;
      RECT 3.64 1.77 3.8 2.855 ;
      RECT 3.64 1.77 5.11 1.935 ;
      RECT 4.84 1.48 5.11 1.935 ;
      RECT 3.865 1.76 5.11 1.935 ;
      RECT 3.865 0.84 4.035 1.935 ;
      RECT 3.59 0.84 4.035 1.09 ;
      RECT 3.14 3.035 4.3 3.205 ;
      RECT 3.99 2.18 4.3 3.205 ;
      RECT 3.14 2.105 3.31 3.205 ;
      RECT 2.11 2.125 2.5 2.415 ;
      RECT 2.33 1.075 2.5 2.415 ;
      RECT 3.3 1.27 3.46 2.27 ;
      RECT 3.3 1.27 3.68 1.59 ;
      RECT 2.33 1.27 3.68 1.435 ;
      RECT 2.11 1.075 2.5 1.35 ;
      RECT 1.52 2.165 1.93 2.355 ;
      RECT 1.77 0.66 1.93 2.355 ;
      RECT 1.77 1.55 2.145 1.88 ;
      RECT 1.455 0.66 1.93 1.25 ;
      RECT 1.455 0.72 3.275 0.89 ;
      RECT 3.105 0.44 3.275 0.89 ;
      RECT 3.105 0.44 4.19 0.63 ;
      RECT 0.38 2.3 0.665 2.945 ;
      RECT 0.38 2.595 2.96 2.755 ;
      RECT 2.79 1.62 2.96 2.755 ;
      RECT 0.38 0.96 0.54 2.945 ;
      RECT 2.79 1.62 3.12 1.92 ;
      RECT 0.38 0.96 0.665 1.27 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhr_1

MACRO sg13g2_dlhrq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhrq_1 0 0 ;
  SIZE 7.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.52 0.6 2 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.185 1.505 1.525 2 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.695 1.57 6.015 2 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6884 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.525 2.075 6.885 3.16 ;
        RECT 6.725 0.77 6.885 3.16 ;
        RECT 6.395 0.77 6.885 1.02 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.2 4 ;
        RECT 6.025 2.205 6.23 4 ;
        RECT 4.875 2.935 5.135 4 ;
        RECT 2.62 2.935 2.88 4 ;
        RECT 0.87 2.935 1.13 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.2 0.22 ;
        RECT 5.905 -0.22 6.165 0.985 ;
        RECT 4.49 -0.22 4.75 0.895 ;
        RECT 2.59 -0.22 2.88 0.745 ;
        RECT 0.995 -0.22 1.26 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.495 2.205 5.735 3.16 ;
      RECT 4.555 2.3 5.735 2.585 ;
      RECT 5.355 1.2 5.515 2.585 ;
      RECT 6.225 1.2 6.545 1.77 ;
      RECT 5.025 1.2 6.545 1.36 ;
      RECT 5.025 0.64 5.285 1.36 ;
      RECT 3.545 2.66 3.785 2.92 ;
      RECT 3.625 1.945 3.785 2.92 ;
      RECT 3.625 1.955 5.175 2.115 ;
      RECT 4.915 1.69 5.175 2.115 ;
      RECT 3.745 0.85 3.905 2.115 ;
      RECT 3.535 0.85 3.905 1.085 ;
      RECT 1.465 2.18 1.875 2.415 ;
      RECT 1.705 1.68 1.875 2.415 ;
      RECT 1.705 1.68 2.08 2 ;
      RECT 4.085 1.445 4.345 1.775 ;
      RECT 1.705 0.925 1.865 2.415 ;
      RECT 4.085 0.475 4.255 1.775 ;
      RECT 1.485 0.605 1.775 1.315 ;
      RECT 1.485 0.925 3.27 1.085 ;
      RECT 3.1 0.475 3.27 1.085 ;
      RECT 3.1 0.475 4.255 0.645 ;
      RECT 3.155 3.18 4.295 3.34 ;
      RECT 3.965 2.295 4.295 3.34 ;
      RECT 3.155 2.195 3.325 3.34 ;
      RECT 2.055 2.2 2.42 2.415 ;
      RECT 2.26 1.265 2.42 2.415 ;
      RECT 3.285 1.265 3.445 2.37 ;
      RECT 3.285 1.265 3.565 1.67 ;
      RECT 2.045 1.265 3.565 1.445 ;
      RECT 0.365 2.37 0.61 3.14 ;
      RECT 0.365 2.595 2.945 2.755 ;
      RECT 2.775 1.69 2.945 2.755 ;
      RECT 0.365 2.37 0.965 2.755 ;
      RECT 0.78 1.12 0.965 2.755 ;
      RECT 2.775 1.69 3.105 2.02 ;
      RECT 0.24 1.12 0.965 1.34 ;
      RECT 0.24 0.92 0.515 1.34 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhrq_1

MACRO sg13g2_dllr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dllr_1 0 0 ;
  SIZE 9.12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 1.48 1.1 2.12 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.29 1.49 1.61 2.12 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.11 1.41 6.45 1.81 ;
    END
  END RESET_B
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.55 2.07 8.96 3.135 ;
        RECT 8.715 0.54 8.96 3.135 ;
        RECT 8.595 0.54 8.96 1.22 ;
    END
  END Q_N
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.245 1.135 7.435 2.2 ;
        RECT 6.89 0.535 7.365 1.25 ;
        RECT 6.975 1.965 7.31 3.035 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 9.12 4 ;
        RECT 8.15 2.06 8.33 4 ;
        RECT 6.455 2.425 6.715 4 ;
        RECT 5.02 2.815 5.695 4 ;
        RECT 2.825 3.12 3.085 4 ;
        RECT 0.905 2.895 1.165 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 9.12 0.22 ;
        RECT 8.085 -0.22 8.345 1.22 ;
        RECT 6.38 -0.22 6.64 1.16 ;
        RECT 5.01 -0.22 5.24 1.165 ;
        RECT 2.785 -0.22 3.045 0.82 ;
        RECT 0.95 -0.22 1.21 1.235 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 7.53 2.355 7.825 2.96 ;
      RECT 7.615 0.725 7.825 2.96 ;
      RECT 7.615 1.52 8.52 1.85 ;
      RECT 7.615 0.725 7.835 1.85 ;
      RECT 7.545 0.725 7.835 0.98 ;
      RECT 5.9 1.99 6.23 3.07 ;
      RECT 4.815 2.2 6.23 2.51 ;
      RECT 6.635 1.48 6.795 2.245 ;
      RECT 5.605 1.99 6.795 2.245 ;
      RECT 5.605 0.555 5.78 2.51 ;
      RECT 6.635 1.48 7.06 1.77 ;
      RECT 5.495 0.555 5.78 1.27 ;
      RECT 3.785 2.625 4.075 2.955 ;
      RECT 3.915 1.855 4.075 2.955 ;
      RECT 3.915 1.855 5.01 2.02 ;
      RECT 4.67 1.44 5.01 2.02 ;
      RECT 4.67 1.44 5.405 1.77 ;
      RECT 4.67 0.595 4.83 2.02 ;
      RECT 3.835 0.595 4.83 0.83 ;
      RECT 3.405 3.155 4.55 3.34 ;
      RECT 4.275 2.27 4.55 3.34 ;
      RECT 3.405 2.2 3.575 3.34 ;
      RECT 1.69 2.43 1.96 2.695 ;
      RECT 1.69 2.43 2.84 2.59 ;
      RECT 2.67 1.35 2.84 2.59 ;
      RECT 1.69 2.41 1.95 2.695 ;
      RECT 1.79 0.595 1.95 2.695 ;
      RECT 3.565 1.35 3.735 2.365 ;
      RECT 2.505 1.465 2.84 1.77 ;
      RECT 3.565 1.35 3.895 1.67 ;
      RECT 2.52 1.35 3.895 1.51 ;
      RECT 1.51 0.595 1.95 1.29 ;
      RECT 2.13 1.955 2.485 2.25 ;
      RECT 2.13 0.605 2.3 2.25 ;
      RECT 4.16 1.01 4.49 1.67 ;
      RECT 2.13 0.605 2.38 1.225 ;
      RECT 2.13 1.01 4.49 1.17 ;
      RECT 2.13 0.605 2.39 1.17 ;
      RECT 1.35 2.95 2.3 3.12 ;
      RECT 2.13 2.78 2.3 3.12 ;
      RECT 0.38 2.355 0.655 3.12 ;
      RECT 1.35 2.355 1.51 3.12 ;
      RECT 2.13 2.78 3.195 2.94 ;
      RECT 3.025 1.69 3.195 2.94 ;
      RECT 0.38 2.355 1.51 2.515 ;
      RECT 0.38 0.875 0.54 3.12 ;
      RECT 3.025 1.69 3.355 2.02 ;
      RECT 0.38 0.875 0.66 1.185 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dllr_1

MACRO sg13g2_dllrq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dllrq_1 0 0 ;
  SIZE 7.68 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.56 1.115 1.96 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.305 1.56 1.62 1.96 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.13 1.29 6.535 1.915 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8449 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.085 2.085 7.415 3.155 ;
        RECT 7.255 0.5 7.415 3.155 ;
        RECT 7.065 0.5 7.415 1.2 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.68 4 ;
        RECT 6.45 2.56 6.705 4 ;
        RECT 4.975 2.7 5.655 4 ;
        RECT 2.715 3.025 2.975 4 ;
        RECT 0.99 2.155 1.25 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.68 0.22 ;
        RECT 6.475 -0.22 6.735 1.105 ;
        RECT 5.01 -0.22 5.27 0.725 ;
        RECT 2.695 -0.22 3.46 0.49 ;
        RECT 0.96 -0.22 1.22 0.49 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.905 2.215 6.165 3.03 ;
      RECT 5.78 0.495 5.95 2.47 ;
      RECT 4.785 2.215 6.885 2.375 ;
      RECT 6.715 1.43 6.885 2.375 ;
      RECT 4.785 2.14 5.95 2.47 ;
      RECT 6.715 1.43 7.075 1.76 ;
      RECT 5.55 0.495 5.95 1.2 ;
      RECT 3.555 2.29 4.035 2.46 ;
      RECT 3.875 1.8 4.035 2.46 ;
      RECT 3.875 1.8 5.37 1.96 ;
      RECT 5.185 1.41 5.37 1.96 ;
      RECT 5.185 1.41 5.595 1.74 ;
      RECT 5.185 0.915 5.355 1.96 ;
      RECT 4.135 0.915 5.355 1.075 ;
      RECT 4.135 0.56 4.395 1.075 ;
      RECT 2.165 2.125 2.545 2.385 ;
      RECT 2.385 1.015 2.545 2.385 ;
      RECT 2.385 1.95 3.69 2.11 ;
      RECT 3.375 1.3 3.69 2.11 ;
      RECT 3.375 1.3 4.635 1.615 ;
      RECT 2.145 1.015 2.545 1.28 ;
      RECT 1.49 2.68 1.975 2.855 ;
      RECT 1.49 2.68 4.545 2.84 ;
      RECT 4.215 2.14 4.545 2.84 ;
      RECT 1.49 2.14 1.965 2.855 ;
      RECT 1.805 1.07 1.965 2.855 ;
      RECT 1.805 1.46 2.205 1.78 ;
      RECT 1.495 1.07 1.965 1.335 ;
      RECT 0.395 2.14 0.75 2.855 ;
      RECT 0.395 0.67 0.565 2.855 ;
      RECT 2.835 0.67 3.165 1.7 ;
      RECT 0.395 0.67 0.745 1.36 ;
      RECT 0.395 0.67 3.165 0.835 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dllrq_1

MACRO sg13g2_dlygate4sd1_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd1_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.24 1.425 0.835 1.945 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.43 2.22 3.685 3.16 ;
        RECT 3.495 0.61 3.685 3.16 ;
        RECT 3.025 1.12 3.685 1.37 ;
        RECT 3.425 0.61 3.685 1.37 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.9 2.455 3.16 4 ;
        RECT 0.91 2.65 1.17 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.915 -0.22 3.175 0.87 ;
        RECT 0.87 -0.22 1.13 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.14 2.03 2.45 2.395 ;
      RECT 2.14 2.03 3.235 2.205 ;
      RECT 3.045 1.55 3.235 2.205 ;
      RECT 2.595 1.55 3.315 1.81 ;
      RECT 2.595 1.16 2.755 1.81 ;
      RECT 2.155 1.16 2.755 1.36 ;
      RECT 2.155 0.96 2.395 1.36 ;
      RECT 1.52 2.615 1.825 2.945 ;
      RECT 1.58 1.57 1.825 2.945 ;
      RECT 1.58 1.57 2.415 1.83 ;
      RECT 1.58 0.615 1.81 2.945 ;
      RECT 1.52 0.615 1.81 0.87 ;
      RECT 0.24 2.195 0.5 2.91 ;
      RECT 0.24 2.195 1.375 2.4 ;
      RECT 1.12 1.065 1.375 2.4 ;
      RECT 0.21 1.065 1.375 1.24 ;
      RECT 0.21 0.61 0.48 1.24 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd1_1

MACRO sg13g2_dlygate4sd2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.425 0.835 1.945 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.43 2.22 3.685 3.16 ;
        RECT 3.495 0.61 3.685 3.16 ;
        RECT 3.065 1.115 3.685 1.37 ;
        RECT 3.425 0.61 3.685 1.37 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.9 2.455 3.16 4 ;
        RECT 0.745 2.65 1.01 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.915 -0.22 3.175 0.87 ;
        RECT 0.86 -0.22 1.12 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.165 2.03 2.425 3.04 ;
      RECT 2.165 2.03 3.205 2.205 ;
      RECT 3.045 1.55 3.205 2.205 ;
      RECT 2.58 1.55 3.315 1.81 ;
      RECT 2.58 1.16 2.74 1.81 ;
      RECT 2.155 1.16 2.74 1.36 ;
      RECT 2.155 0.96 2.395 1.36 ;
      RECT 1.52 2.615 1.825 2.945 ;
      RECT 1.58 1.555 1.825 2.945 ;
      RECT 1.58 1.555 2.4 1.815 ;
      RECT 1.58 0.61 1.81 2.945 ;
      RECT 1.52 0.61 1.81 0.87 ;
      RECT 0.24 2.195 0.5 2.91 ;
      RECT 0.24 2.195 1.375 2.4 ;
      RECT 1.12 1.065 1.375 2.4 ;
      RECT 0.21 1.065 1.375 1.24 ;
      RECT 0.21 0.61 0.48 1.24 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd2_1

MACRO sg13g2_dlygate4sd3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd3_1 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1.41 0.915 2.08 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.12 2.56 3.38 4 ;
        RECT 0.81 2.665 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.13 -0.22 3.39 0.85 ;
        RECT 0.8 -0.22 1.07 0.835 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 2.075 4.02 3.17 ;
        RECT 3.805 0.595 4.02 3.17 ;
        RECT 3.61 0.595 4.02 1.34 ;
    END
  END X
  OBS
    LAYER Metal1 ;
      RECT 2.21 2.045 2.47 3.04 ;
      RECT 2.21 2.045 3.34 2.215 ;
      RECT 3.15 1.045 3.34 2.215 ;
      RECT 3.15 1.515 3.535 1.845 ;
      RECT 2.205 1.045 3.34 1.235 ;
      RECT 2.205 0.945 2.47 1.235 ;
      RECT 1.69 2.22 1.955 3.16 ;
      RECT 1.72 0.665 1.955 3.16 ;
      RECT 1.72 1.55 2.925 1.81 ;
      RECT 0.3 2.32 0.56 2.88 ;
      RECT 0.3 2.32 1.455 2.48 ;
      RECT 1.175 1.015 1.455 2.48 ;
      RECT 0.3 1.015 1.455 1.205 ;
      RECT 0.3 0.69 0.56 1.205 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd3_1

MACRO sg13g2_ebufn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_2 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5044 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 1.37 3.495 1.85 ;
    END
  END TE_B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.695 1.37 4.015 1.85 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 2.17 1.1 2.765 ;
        RECT 0.74 0.845 1.025 1.08 ;
        RECT 0.74 0.845 0.91 2.38 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 3.52 2.915 3.78 4 ;
        RECT 1.89 3.23 2.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 3.56 -0.22 3.82 1.13 ;
        RECT 1.78 -0.22 2.04 0.82 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 4.14 2.08 4.435 3.04 ;
      RECT 4.245 0.595 4.435 3.04 ;
      RECT 2.36 2.545 4.435 2.71 ;
      RECT 2.36 1.6 2.52 2.71 ;
      RECT 1.1 1.6 2.52 1.76 ;
      RECT 1.1 1.5 1.355 1.76 ;
      RECT 4.06 0.595 4.435 1.13 ;
      RECT 2.7 2.08 3.22 2.34 ;
      RECT 2.7 0.975 2.915 2.34 ;
      RECT 2.7 0.975 3.3 1.16 ;
      RECT 3.05 0.56 3.3 1.16 ;
      RECT 0.33 3.075 1.61 3.235 ;
      RECT 1.35 2.17 1.61 3.235 ;
      RECT 2.43 2.89 2.69 3.16 ;
      RECT 0.33 2.51 0.59 3.235 ;
      RECT 1.35 2.89 2.69 3.05 ;
      RECT 1.27 1 2.515 1.16 ;
      RECT 2.3 0.54 2.515 1.16 ;
      RECT 0.25 0.44 0.51 1.16 ;
      RECT 1.27 0.44 1.53 1.16 ;
      RECT 0.25 0.44 1.53 0.635 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_2

MACRO sg13g2_ebufn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_4 0 0 ;
  SIZE 7.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.96 1.185 2.24 ;
        RECT 0.65 1.535 0.915 2.24 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8242 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 1.42 1.855 1.7 ;
        RECT 1.3 1.02 1.58 1.7 ;
    END
  END TE_B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4322 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.15 2.11 6.41 2.83 ;
        RECT 6.23 0.93 6.41 2.83 ;
        RECT 5.115 1.145 6.41 1.375 ;
        RECT 6.145 0.93 6.41 1.375 ;
        RECT 5.12 2.11 6.41 2.335 ;
        RECT 5.12 2.11 5.38 2.83 ;
        RECT 5.115 0.93 5.375 1.375 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.2 4 ;
        RECT 4.09 2.57 4.35 4 ;
        RECT 3.07 2.945 3.33 4 ;
        RECT 0.89 2.91 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.2 0.22 ;
        RECT 4.09 -0.22 4.35 1.16 ;
        RECT 3.07 -0.22 3.33 1.16 ;
        RECT 0.805 -0.22 1.065 1.19 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.56 1.34 4.82 1.51 ;
      RECT 4.6 0.455 4.82 1.51 ;
      RECT 3.58 0.59 3.84 1.51 ;
      RECT 2.56 0.59 2.82 1.51 ;
      RECT 6.66 0.455 6.92 1.19 ;
      RECT 5.635 0.455 5.895 0.85 ;
      RECT 4.6 0.455 6.92 0.625 ;
      RECT 4.615 3.17 6.92 3.33 ;
      RECT 6.66 2.23 6.92 3.33 ;
      RECT 3.58 2.115 3.84 3.17 ;
      RECT 2.56 2.6 2.82 3.17 ;
      RECT 5.64 2.57 5.9 3.33 ;
      RECT 4.615 2.115 4.845 3.33 ;
      RECT 2.56 2.6 3.84 2.765 ;
      RECT 3.58 2.115 4.845 2.275 ;
      RECT 0.28 2.555 0.64 3.17 ;
      RECT 0.28 2.57 2.12 2.73 ;
      RECT 1.96 2.23 2.12 2.73 ;
      RECT 0.28 0.59 0.445 3.17 ;
      RECT 1.96 2.23 3.2 2.39 ;
      RECT 3.03 1.7 3.2 2.39 ;
      RECT 3.03 1.7 5.935 1.86 ;
      RECT 4.995 1.595 5.935 1.86 ;
      RECT 0.28 0.59 0.54 1.19 ;
      RECT 1.4 1.885 1.66 2.39 ;
      RECT 1.4 1.885 2.355 2.05 ;
      RECT 2.095 0.535 2.355 2.05 ;
      RECT 1.315 0.59 2.355 0.84 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_4

MACRO sg13g2_ebufn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_8 0 0 ;
  SIZE 12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.73 2.12 3.99 2.85 ;
        RECT 0.67 1.17 3.99 1.36 ;
        RECT 3.73 0.915 3.99 1.36 ;
        RECT 0.67 2.12 3.99 2.29 ;
        RECT 2.71 2.12 2.97 2.85 ;
        RECT 2.71 0.92 2.97 1.36 ;
        RECT 0.67 2.12 2.97 2.295 ;
        RECT 1.69 2.12 1.95 2.85 ;
        RECT 1.685 0.92 1.95 1.36 ;
        RECT 0.78 1.17 1.14 2.295 ;
        RECT 0.67 2.02 0.93 2.85 ;
        RECT 0.67 0.92 0.93 1.465 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.84 1.51 11.335 1.835 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.665 1.51 10.605 1.835 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12 4 ;
        RECT 11.51 2.62 11.77 4 ;
        RECT 10.49 2.93 10.75 4 ;
        RECT 7.84 3.205 8.105 4 ;
        RECT 6.795 2.96 7.055 4 ;
        RECT 5.77 2.96 6.03 4 ;
        RECT 4.75 2.97 5.01 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12 0.22 ;
        RECT 11.51 -0.22 11.77 0.9 ;
        RECT 10.49 -0.22 10.75 1.24 ;
        RECT 7.875 -0.22 8.135 1.225 ;
        RECT 6.855 -0.22 7.115 1.225 ;
        RECT 5.835 -0.22 6.095 1.225 ;
        RECT 4.815 -0.22 5.075 1.2 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 11 2.24 11.26 3.19 ;
      RECT 8.805 2.56 11.26 2.725 ;
      RECT 8.805 2.25 8.985 2.725 ;
      RECT 11 2.24 11.765 2.44 ;
      RECT 11.59 1.08 11.765 2.44 ;
      RECT 4.235 2.25 8.985 2.41 ;
      RECT 4.235 1.73 4.445 2.41 ;
      RECT 1.58 1.73 4.445 1.9 ;
      RECT 1.58 1.585 3.995 1.9 ;
      RECT 11 1.08 11.765 1.24 ;
      RECT 11 0.64 11.26 1.24 ;
      RECT 9.165 2.1 10.24 2.38 ;
      RECT 9.165 0.64 9.4 2.38 ;
      RECT 9.98 0.64 10.24 1.24 ;
      RECT 8.875 0.64 10.24 0.885 ;
      RECT 4.72 1.55 8.645 1.72 ;
      RECT 8.385 0.74 8.645 1.72 ;
      RECT 4.26 1.38 5.585 1.55 ;
      RECT 7.365 0.74 7.625 1.72 ;
      RECT 6.345 0.74 6.605 1.72 ;
      RECT 5.325 0.74 5.585 1.72 ;
      RECT 4.26 0.53 4.525 1.55 ;
      RECT 0.15 0.53 0.405 1.34 ;
      RECT 3.22 0.53 3.48 0.985 ;
      RECT 2.2 0.53 2.46 0.985 ;
      RECT 1.18 0.53 1.44 0.975 ;
      RECT 0.15 0.53 4.525 0.73 ;
      RECT 0.16 3.155 4.5 3.325 ;
      RECT 4.24 2.59 4.5 3.325 ;
      RECT 8.385 2.84 8.645 3.19 ;
      RECT 7.305 2.59 7.565 3.19 ;
      RECT 6.285 2.59 6.55 3.19 ;
      RECT 5.26 2.59 5.52 3.19 ;
      RECT 3.22 2.59 3.48 3.325 ;
      RECT 2.2 2.59 2.46 3.325 ;
      RECT 1.18 2.59 1.44 3.325 ;
      RECT 0.16 2.15 0.42 3.325 ;
      RECT 7.305 2.84 8.645 3.02 ;
      RECT 4.24 2.59 6.55 2.78 ;
      RECT 4.24 2.59 7.565 2.775 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_8

MACRO sg13g2_einvn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7142 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.16 1.005 3.49 2.825 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.7 1.01 4.03 1.75 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.429 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 1.32 0.995 2.33 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 2.14 2.56 2.4 4 ;
        RECT 0.6 2.56 0.86 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 2.14 -0.22 2.4 0.85 ;
        RECT 0.6 -0.22 0.865 0.91 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.655 1.03 2.91 1.195 ;
      RECT 2.65 0.59 2.91 1.195 ;
      RECT 1.655 0.575 1.9 1.195 ;
      RECT 2.65 0.59 3.95 0.825 ;
      RECT 2.65 3.175 3.93 3.335 ;
      RECT 3.67 2.22 3.93 3.335 ;
      RECT 2.65 2.215 2.91 3.335 ;
      RECT 1.63 2.215 1.89 3.16 ;
      RECT 1.63 2.215 2.91 2.38 ;
      RECT 1.085 2.56 1.385 3.16 ;
      RECT 1.215 1.52 1.385 3.16 ;
      RECT 1.215 1.52 1.655 1.85 ;
      RECT 1.215 0.65 1.38 3.16 ;
      RECT 1.115 0.65 1.38 0.91 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_2

MACRO sg13g2_einvn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_4 0 0 ;
  SIZE 6.24 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.2 1.115 5.56 1.305 ;
        RECT 5.3 0.89 5.56 1.305 ;
        RECT 5.1 2.13 5.36 2.82 ;
        RECT 4.08 2.13 5.36 2.33 ;
        RECT 4.2 1.025 4.54 1.305 ;
        RECT 4.2 1.025 4.435 2.33 ;
        RECT 4.08 2.015 4.34 2.82 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.65 1.54 5.59 1.925 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8242 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 1.46 0.725 2 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 6.24 4 ;
        RECT 3.06 2.22 3.32 4 ;
        RECT 2.04 2.22 2.3 4 ;
        RECT 0.365 2.22 0.625 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 6.24 0.22 ;
        RECT 3.26 -0.22 3.52 1.21 ;
        RECT 2.24 -0.22 2.5 1.21 ;
        RECT 0.365 -0.22 0.625 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.77 1.405 4 1.575 ;
      RECT 3.77 0.605 4 1.575 ;
      RECT 2.75 0.61 3.01 1.575 ;
      RECT 1.77 0.61 1.965 1.575 ;
      RECT 5.81 0.475 6.07 1.21 ;
      RECT 3.77 0.605 5.06 0.84 ;
      RECT 4.77 0.475 6.07 0.645 ;
      RECT 3.57 3.14 5.87 3.335 ;
      RECT 5.61 2.22 5.87 3.335 ;
      RECT 2.55 1.795 2.81 3.16 ;
      RECT 1.53 1.795 1.79 3.16 ;
      RECT 4.59 2.54 4.85 3.335 ;
      RECT 3.57 1.795 3.83 3.335 ;
      RECT 1.53 1.795 3.83 2.01 ;
      RECT 0.875 2.22 1.135 3.16 ;
      RECT 0.91 0.61 1.135 3.16 ;
      RECT 0.875 0.61 1.57 1.21 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_4

MACRO sg13g2_einvn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_8 0 0 ;
  SIZE 10.56 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.9344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.43 1.51 9.84 1.845 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.33 2.12 9.59 2.815 ;
        RECT 6.26 1.09 9.59 1.28 ;
        RECT 9.33 0.915 9.59 1.28 ;
        RECT 6.26 2.12 9.59 2.31 ;
        RECT 8.31 2.12 8.57 2.815 ;
        RECT 8.31 0.925 8.57 1.28 ;
        RECT 7.29 2.12 7.55 2.815 ;
        RECT 7.29 1.055 7.55 1.28 ;
        RECT 6.26 1.09 6.955 2.31 ;
        RECT 6.26 1.055 6.525 2.77 ;
    END
  END Z
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.37 0.63 1.82 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 10.56 4 ;
        RECT 4.985 2.565 5.245 4 ;
        RECT 3.965 2.245 4.225 4 ;
        RECT 2.945 2.245 3.205 4 ;
        RECT 1.925 2.245 2.185 4 ;
        RECT 0.35 2.08 0.61 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 10.56 0.22 ;
        RECT 5.25 -0.22 5.51 1.21 ;
        RECT 4.23 -0.22 4.49 1.3 ;
        RECT 3.21 -0.22 3.47 1.3 ;
        RECT 2.19 -0.22 2.45 1.3 ;
        RECT 0.355 -0.22 0.615 1.18 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.72 1.49 6.005 1.66 ;
      RECT 5.765 0.57 6.005 1.66 ;
      RECT 4.74 0.665 5 1.66 ;
      RECT 3.72 0.67 3.98 1.66 ;
      RECT 2.7 0.67 2.96 1.66 ;
      RECT 1.72 0.615 1.93 1.66 ;
      RECT 9.84 0.445 10.1 1.305 ;
      RECT 8.82 0.445 9.08 0.9 ;
      RECT 7.8 0.445 8.06 0.885 ;
      RECT 6.78 0.57 7.04 0.855 ;
      RECT 5.765 0.57 8.06 0.79 ;
      RECT 7.795 0.445 10.1 0.615 ;
      RECT 5.75 3.085 10.1 3.295 ;
      RECT 9.84 2.245 10.1 3.295 ;
      RECT 1.41 1.885 1.67 3.13 ;
      RECT 4.475 2.17 4.735 3.12 ;
      RECT 3.455 1.885 3.715 3.12 ;
      RECT 2.435 1.885 2.695 3.12 ;
      RECT 8.82 2.575 9.08 3.295 ;
      RECT 7.8 2.55 8.06 3.295 ;
      RECT 6.78 2.58 7.045 3.295 ;
      RECT 5.75 2.17 6.025 3.295 ;
      RECT 4.475 2.17 6.025 2.34 ;
      RECT 4.475 1.885 4.69 3.12 ;
      RECT 1.41 1.885 4.69 2.055 ;
      RECT 0.86 1.32 1.12 3.13 ;
      RECT 0.88 0.575 1.52 1.525 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_8

MACRO sg13g2_fill_1
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_1 0 0 ;
  SIZE 0.48 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 0.48 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 0.48 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_1

MACRO sg13g2_fill_2
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_2 0 0 ;
  SIZE 0.96 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 0.96 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 0.96 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_2

MACRO sg13g2_fill_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_4 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_4

MACRO sg13g2_fill_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_8 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_8

MACRO sg13g2_inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_1 0 0 ;
  SIZE 1.44 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.44 4 ;
        RECT 0.33 2.235 0.59 4 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.855 0.61 1.085 3.175 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 1.52 0.625 1.85 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.44 0.22 ;
        RECT 0.33 -0.22 0.59 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_1

MACRO sg13g2_inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_16 0 0 ;
  SIZE 9.12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 3.8688 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.025 1.49 8.785 1.87 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.6544 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.975 2.145 8.235 3.16 ;
        RECT 6.955 1.05 8.235 1.21 ;
        RECT 7.975 0.625 8.235 1.21 ;
        RECT 0.835 2.145 8.235 2.32 ;
        RECT 6.955 0.625 7.215 3.16 ;
        RECT 0.835 1.9 7.215 2.32 ;
        RECT 5.935 0.625 6.195 3.16 ;
        RECT 4.915 0.625 5.175 3.16 ;
        RECT 3.895 0.625 4.155 3.16 ;
        RECT 2.875 0.625 3.135 3.16 ;
        RECT 1.855 0.63 2.115 3.16 ;
        RECT 0.835 0.63 1.095 3.16 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 9.12 4 ;
        RECT 7.465 3.555 8.795 4 ;
        RECT 8.535 2.22 8.795 4 ;
        RECT 7.465 2.56 7.725 4 ;
        RECT 6.445 2.56 6.705 4 ;
        RECT 5.425 2.56 5.685 4 ;
        RECT 4.405 2.56 4.665 4 ;
        RECT 3.385 2.56 3.645 4 ;
        RECT 2.365 2.56 2.625 4 ;
        RECT 1.345 2.56 1.605 4 ;
        RECT 0.325 2.22 0.585 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 9.12 0.22 ;
        RECT 8.485 -0.22 8.745 1.21 ;
        RECT 7.465 -0.22 7.725 0.87 ;
        RECT 6.445 -0.22 6.705 1.21 ;
        RECT 5.425 -0.22 5.685 1.21 ;
        RECT 4.405 -0.22 4.665 1.21 ;
        RECT 3.385 -0.22 3.645 1.21 ;
        RECT 2.365 -0.22 2.625 1.21 ;
        RECT 1.345 -0.22 1.605 1.21 ;
        RECT 0.325 -0.22 0.585 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_16

MACRO sg13g2_inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_2 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 1.52 1.59 1.85 ;
        RECT 0.795 2.22 1.055 3.18 ;
        RECT 0.87 0.61 1.055 3.18 ;
        RECT 0.795 0.61 1.055 1.21 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1.52 0.635 1.85 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.31 2.22 1.57 4 ;
        RECT 0.285 2.22 0.545 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.305 -0.22 1.565 1.21 ;
        RECT 0.285 -0.22 0.545 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_2

MACRO sg13g2_inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_4 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 1.52 2 1.9 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 2.17 2.54 2.34 ;
        RECT 2.245 1.05 2.54 2.34 ;
        RECT 0.775 1.05 2.54 1.21 ;
        RECT 1.795 2.17 2.055 3.155 ;
        RECT 1.795 0.61 2.055 1.21 ;
        RECT 0.775 2.17 1.035 3.155 ;
        RECT 0.775 0.61 1.035 1.21 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.305 2.545 2.565 4 ;
        RECT 1.285 2.545 1.545 4 ;
        RECT 0.265 2.205 0.525 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.305 -0.22 2.565 0.87 ;
        RECT 1.28 -0.22 1.55 0.87 ;
        RECT 0.265 -0.22 0.525 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_4

MACRO sg13g2_inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_8 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8458 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.775 0.61 4.035 3.16 ;
        RECT 2.74 1.53 4.035 1.84 ;
        RECT 2.755 0.61 3.015 3.16 ;
        RECT 0.715 2.22 3.015 2.38 ;
        RECT 2.74 1.07 3.015 2.38 ;
        RECT 0.715 1.07 3.015 1.23 ;
        RECT 0.715 1.05 2 1.23 ;
        RECT 1.735 0.61 2 1.23 ;
        RECT 1.735 2.22 1.995 3.16 ;
        RECT 0.715 0.62 0.98 1.23 ;
        RECT 0.715 2.22 0.975 3.16 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.9344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 1.535 2.495 1.865 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 4.295 2.22 4.555 4 ;
        RECT 3.265 2.22 3.525 4 ;
        RECT 2.245 2.56 2.505 4 ;
        RECT 1.225 2.56 1.485 4 ;
        RECT 0.205 2.22 0.465 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 4.295 -0.22 4.555 1.21 ;
        RECT 3.265 -0.22 3.525 1.21 ;
        RECT 2.245 -0.22 2.505 0.89 ;
        RECT 1.225 -0.22 1.485 0.87 ;
        RECT 0.205 -0.22 0.465 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_8

MACRO sg13g2_lgcp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_lgcp_1 0 0 ;
  SIZE 7.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.68 1.635 2.21 ;
    END
  END GATE
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3978 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.68 1.685 5.125 2.015 ;
        RECT 4.68 1.685 4.955 2.42 ;
    END
  END CLK
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.495 1.76 6.845 3.16 ;
        RECT 6.59 0.56 6.845 3.16 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.2 4 ;
        RECT 5.99 2.2 6.25 4 ;
        RECT 4.72 2.73 4.98 4 ;
        RECT 3.115 3.095 3.38 4 ;
        RECT 0.89 2.89 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.2 0.22 ;
        RECT 6.09 -0.22 6.35 1.26 ;
        RECT 4.69 -0.22 4.95 1.445 ;
        RECT 2.99 0.895 3.525 1.125 ;
        RECT 3.365 -0.22 3.525 1.125 ;
        RECT 0.9 -0.22 1.115 0.8 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.23 2.195 5.49 2.995 ;
      RECT 5.23 2.195 5.765 2.355 ;
      RECT 5.585 0.815 5.765 2.355 ;
      RECT 5.585 1.51 6.275 1.84 ;
      RECT 5.585 0.815 5.855 1.84 ;
      RECT 5.525 0.815 5.855 1.41 ;
      RECT 4.205 2.155 4.47 2.995 ;
      RECT 3.115 2.695 4.47 2.905 ;
      RECT 3.115 1.725 3.29 2.905 ;
      RECT 1.975 2.305 3.29 2.565 ;
      RECT 1.975 1.36 2.235 2.565 ;
      RECT 4.205 1.23 4.445 2.995 ;
      RECT 3.115 1.725 3.655 2.04 ;
      RECT 3.65 2.26 4.015 2.45 ;
      RECT 3.845 0.845 4.015 2.45 ;
      RECT 2.445 1.37 2.775 2.05 ;
      RECT 2.445 1.37 4.015 1.54 ;
      RECT 3.705 0.845 4.015 1.54 ;
      RECT 0.35 2.125 0.61 3.15 ;
      RECT 0.33 1.05 0.495 2.48 ;
      RECT 0.35 0.6 0.595 1.3 ;
      RECT 1.295 0.465 1.455 1.16 ;
      RECT 0.35 0.98 1.455 1.16 ;
      RECT 2.865 0.465 3.185 0.71 ;
      RECT 1.295 0.465 3.185 0.635 ;
      RECT 1.625 2.795 2.35 3.055 ;
      RECT 1.625 2.42 1.785 3.055 ;
      RECT 0.855 2.42 1.785 2.58 ;
      RECT 0.855 1.34 1.025 2.58 ;
      RECT 0.675 1.51 1.025 1.84 ;
      RECT 0.855 1.34 1.795 1.5 ;
      RECT 1.635 0.89 1.795 1.5 ;
      RECT 1.635 0.89 2.395 1.14 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_lgcp_1

MACRO sg13g2_mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux2_1 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.4 2.535 1.92 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.92 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.5 1.105 1.87 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0081 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.135 2.04 4.59 3.2 ;
        RECT 4.4 0.57 4.59 3.2 ;
        RECT 4.315 0.57 4.59 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.855 2.345 2.56 2.505 ;
      RECT 1.855 2.08 2.015 2.505 ;
      RECT 1.285 2.08 2.015 2.26 ;
      RECT 1.285 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.22 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.285 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.295 2.28 0.575 2.88 ;
      RECT 0.295 2.44 1.64 2.6 ;
      RECT 0.295 0.8 0.455 2.88 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.295 0.8 0.575 1.06 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux2_1

MACRO sg13g2_mux2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux2_2 0 0 ;
  SIZE 5.28 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.175 1.4 2.535 1.875 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.785 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.5 1.11 1.905 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.023 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.135 2.04 4.685 3.2 ;
        RECT 4.515 0.61 4.685 3.2 ;
        RECT 4.315 0.61 4.685 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 5.28 4 ;
        RECT 4.905 2.08 5.105 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 5.28 0.22 ;
        RECT 4.875 -0.22 5.135 1.21 ;
        RECT 3.6 -0.22 3.86 0.87 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.825 2.345 2.56 2.505 ;
      RECT 1.825 2.1 1.985 2.505 ;
      RECT 1.29 2.1 1.985 2.26 ;
      RECT 1.29 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.245 1.85 ;
      RECT 3.945 1.1 4.135 1.85 ;
      RECT 3.195 1.1 4.135 1.26 ;
      RECT 3.195 0.61 3.365 1.26 ;
      RECT 1.29 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.45 3.295 ;
      RECT 3.29 1.54 3.45 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.31 2.28 0.575 2.88 ;
      RECT 0.31 2.44 1.64 2.6 ;
      RECT 0.31 0.92 0.47 2.88 ;
      RECT 3.29 1.54 3.72 1.87 ;
      RECT 0.31 0.92 0.575 1.18 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux2_2

MACRO sg13g2_mux4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux4_1 0 0 ;
  SIZE 10.08 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6396 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 1.435 1.095 1.92 ;
    END
  END S0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 1.435 1.57 1.92 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.22 1.435 3.54 2.255 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.72 1.435 4.09 2.255 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.07 1.53 6.4 1.96 ;
    END
  END A3
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4264 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.52 1.56 8.955 1.895 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.64 2.78 9.905 3.075 ;
        RECT 9.665 0.62 9.905 3.075 ;
        RECT 9.475 0.62 9.905 1.36 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 10.08 4 ;
        RECT 9.095 2.585 9.355 4 ;
        RECT 5.95 2.905 6.28 4 ;
        RECT 3.52 2.92 3.78 4 ;
        RECT 0.985 2.12 1.245 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 10.08 0.22 ;
        RECT 9.035 -0.22 9.295 1.325 ;
        RECT 5.545 -0.22 5.805 0.96 ;
        RECT 3.495 -0.22 3.77 0.835 ;
        RECT 0.985 -0.22 1.245 0.84 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 7.01 3.125 8.91 3.295 ;
      RECT 8.75 2.23 8.91 3.295 ;
      RECT 7.01 1.335 7.3 3.295 ;
      RECT 8.75 2.23 9.46 2.4 ;
      RECT 9.2 1.605 9.46 2.4 ;
      RECT 6.965 1.16 7.21 1.505 ;
      RECT 8.195 2.205 8.57 2.81 ;
      RECT 8.195 1.97 8.355 2.81 ;
      RECT 8.17 1.97 8.355 2.2 ;
      RECT 8.18 1.4 8.34 2.2 ;
      RECT 7.85 1.665 8.34 1.995 ;
      RECT 8.195 0.76 8.355 1.485 ;
      RECT 8.195 0.76 8.745 1.36 ;
      RECT 4.525 2.2 5.385 2.945 ;
      RECT 7.51 2.22 7.86 2.81 ;
      RECT 4.525 2.2 5.885 2.37 ;
      RECT 5.715 1.14 5.885 2.37 ;
      RECT 7.51 1.26 7.67 2.81 ;
      RECT 7.51 1.26 7.98 1.42 ;
      RECT 7.845 0.44 8.005 1.35 ;
      RECT 5.15 1.14 6.375 1.3 ;
      RECT 6.115 0.44 6.375 1.3 ;
      RECT 5.15 0.595 5.32 1.3 ;
      RECT 4.55 0.595 5.32 0.87 ;
      RECT 6.115 0.44 8.005 0.6 ;
      RECT 4.015 3.125 5.77 3.295 ;
      RECT 5.57 2.555 5.77 3.295 ;
      RECT 6.51 2.17 6.78 3.16 ;
      RECT 6.58 0.82 6.78 3.16 ;
      RECT 4.015 2.435 4.24 3.295 ;
      RECT 2.26 1.95 2.77 2.905 ;
      RECT 5.57 2.555 6.78 2.725 ;
      RECT 2.26 2.435 4.24 2.595 ;
      RECT 2.26 0.87 2.42 2.905 ;
      RECT 2.095 0.87 2.42 1.2 ;
      RECT 7.45 0.82 7.665 1.08 ;
      RECT 6.58 0.82 7.665 0.98 ;
      RECT 0.33 2.12 0.745 2.985 ;
      RECT 0.33 0.59 0.5 2.985 ;
      RECT 4.8 1.665 5.535 1.97 ;
      RECT 1.75 1.42 2.08 1.75 ;
      RECT 4.3 1.05 4.61 1.67 ;
      RECT 2.68 1.05 3.01 1.67 ;
      RECT 4.8 1.05 4.97 1.97 ;
      RECT 1.75 0.475 1.915 1.75 ;
      RECT 2.68 1.05 4.97 1.21 ;
      RECT 0.33 1.02 1.915 1.2 ;
      RECT 2.68 0.475 2.85 1.67 ;
      RECT 0.33 0.59 0.64 1.2 ;
      RECT 1.75 0.475 2.85 0.645 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux4_1

MACRO sg13g2_nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.83 1.06 1.6 1.245 ;
        RECT 1.34 0.62 1.6 1.245 ;
        RECT 0.83 1.06 1.09 3.16 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.27 1.47 1.6 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 1.47 0.62 1.9 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.34 2.08 1.6 4 ;
        RECT 0.32 2.08 0.58 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.32 -0.22 0.58 1.275 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2_1

MACRO sg13g2_nand2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1248 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.88 2.5 2.14 3.16 ;
        RECT 1.32 1.39 2.14 1.55 ;
        RECT 1.88 1 2.14 1.55 ;
        RECT 0.85 2.5 2.14 2.72 ;
        RECT 1.32 1.39 1.56 2.72 ;
        RECT 0.85 2.5 1.11 3.16 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 1.73 2.17 1.98 ;
        RECT 1.79 1.73 2.05 2.32 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.435 1.1 1.9 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.39 2.16 2.65 4 ;
        RECT 1.36 2.9 1.62 4 ;
        RECT 0.32 2.08 0.58 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 0.85 -0.22 1.11 0.855 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.37 0.53 2.65 1.2 ;
      RECT 0.325 1.035 1.62 1.2 ;
      RECT 1.35 0.53 1.62 1.2 ;
      RECT 0.325 0.5 0.585 1.2 ;
      RECT 1.35 0.53 2.65 0.76 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2_2

MACRO sg13g2_nand2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2b_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7586 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 2.54 2.16 2.7 ;
        RECT 2 0.61 2.16 2.7 ;
        RECT 1.745 0.61 2.16 1.315 ;
        RECT 1.205 2.54 1.465 3.16 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.53 1.205 1.835 ;
    END
  END B
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 1.53 0.6 1.835 ;
    END
  END A_N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.715 2.9 1.975 4 ;
        RECT 0.695 2.54 0.955 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.69 -0.22 0.96 0.94 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.155 2.17 0.415 2.88 ;
      RECT 0.155 2.17 1.545 2.355 ;
      RECT 1.385 1.19 1.545 2.355 ;
      RECT 1.385 1.52 1.805 1.83 ;
      RECT 0.155 1.19 1.545 1.35 ;
      RECT 0.155 0.92 0.415 1.35 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2b_1

MACRO sg13g2_nand2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2b_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1248 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.71 2.2 3 3.18 ;
        RECT 2.77 1 3 3.18 ;
        RECT 2.71 1 3 1.39 ;
        RECT 1.68 2.2 3 2.36 ;
        RECT 1.68 2.2 1.94 3.16 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.16 1.535 2.59 1.845 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.22 2.22 3.48 4 ;
        RECT 2.19 2.56 2.45 4 ;
        RECT 1.15 2.125 1.41 4 ;
        RECT 0.13 2.28 0.39 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 1.68 -0.22 1.94 0.855 ;
        RECT 0.13 -0.22 0.39 1.275 ;
    END
  END VSS
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.155 1.475 0.61 1.865 ;
    END
  END A_N
  OBS
    LAYER Metal1 ;
      RECT 3.2 0.53 3.48 1.2 ;
      RECT 1.155 1.035 2.45 1.2 ;
      RECT 2.18 0.53 2.45 1.2 ;
      RECT 1.155 0.6 1.415 1.2 ;
      RECT 2.18 0.53 3.48 0.76 ;
      RECT 0.64 2.21 0.9 2.88 ;
      RECT 0.805 1.015 0.965 2.34 ;
      RECT 0.805 1.585 1.47 1.845 ;
      RECT 0.64 1.015 0.965 1.275 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2b_2

MACRO sg13g2_nand3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand3_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.505 1.22 1.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.505 0.65 1.89 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.745 1.505 2.155 1.89 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.058 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 2.29 2.07 3.23 ;
        RECT 1.4 0.975 2.07 1.23 ;
        RECT 1.81 0.63 2.07 1.23 ;
        RECT 0.79 2.29 2.07 2.45 ;
        RECT 1.4 0.975 1.565 2.45 ;
        RECT 0.79 2.29 1.05 3.23 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.3 2.63 1.56 4 ;
        RECT 0.28 2.29 0.54 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.28 -0.22 0.54 1.23 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand3_1

MACRO sg13g2_nand3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand3b_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 1.475 2.1 1.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 1.475 1.62 1.9 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1468 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.67 2.2 3.13 3.16 ;
        RECT 2.96 0.63 3.13 3.16 ;
        RECT 2.775 0.63 3.13 1.23 ;
        RECT 1.65 2.2 3.13 2.39 ;
        RECT 1.65 2.2 1.91 3.16 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.16 2.575 2.42 4 ;
        RECT 1.14 2.22 1.4 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 1.08 -0.22 1.35 0.89 ;
    END
  END VSS
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 1.475 1.08 1.9 ;
    END
  END A_N
  OBS
    LAYER Metal1 ;
      RECT 0.44 2.28 0.86 2.88 ;
      RECT 0.44 0.945 0.61 2.88 ;
      RECT 2.43 1.59 2.755 1.85 ;
      RECT 2.43 1.07 2.59 1.85 ;
      RECT 0.44 1.07 2.59 1.23 ;
      RECT 0.44 0.945 0.75 1.23 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand3b_1

MACRO sg13g2_nand4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand4_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 1.59 1.7 1.85 ;
        RECT 1.44 1.14 1.64 1.85 ;
        RECT 1.32 1.14 1.64 1.38 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.55 1.19 1.87 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.965 1.59 2.24 1.85 ;
        RECT 1.965 1.27 2.125 1.85 ;
        RECT 1.8 0.72 2.04 0.96 ;
        RECT 1.84 0.72 2 1.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1028 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 2.29 2.62 2.45 ;
        RECT 2.46 0.63 2.62 2.45 ;
        RECT 2.32 0.63 2.62 1.23 ;
        RECT 1.8 2.29 2.07 3.225 ;
        RECT 0.79 2.29 1.05 3.225 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.32 2.63 2.58 4 ;
        RECT 1.3 2.63 1.56 4 ;
        RECT 0.28 2.29 0.54 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 0.28 -0.22 0.54 1.23 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.55 0.6 1.87 ;
    END
  END D
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand4_1

MACRO sg13g2_nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.35 1.52 0.68 1.85 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.52 1.58 1.85 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 2.235 1.57 3.16 ;
        RECT 0.87 2.235 1.57 2.435 ;
        RECT 0.87 0.605 1.17 1.21 ;
        RECT 0.87 0.605 1.04 2.435 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.4 2.22 0.66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.42 -0.22 1.68 1.21 ;
        RECT 0.4 -0.22 0.66 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2_1

MACRO sg13g2_nor2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.53 1.13 1.84 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.77 1.53 2.15 1.84 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.988 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 2.22 2.6 2.38 ;
        RECT 2.44 1.075 2.6 2.38 ;
        RECT 0.81 1.075 2.6 1.24 ;
        RECT 1.78 2.22 2.09 2.72 ;
        RECT 1.83 0.59 2.085 1.24 ;
        RECT 0.81 0.61 1.065 1.24 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 0.81 2.56 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.34 -0.22 2.6 0.865 ;
        RECT 1.32 -0.22 1.58 0.87 ;
        RECT 0.3 -0.22 0.56 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.32 2.9 2.6 3.16 ;
      RECT 2.34 2.56 2.6 3.16 ;
      RECT 0.3 2.22 0.56 3.16 ;
      RECT 1.32 2.22 1.58 3.16 ;
      RECT 0.3 2.22 1.58 2.38 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2_2

MACRO sg13g2_nor2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2b_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 1.5 2.06 1.87 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.27 1.5 0.62 1.87 ;
    END
  END B_N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 2.235 2.06 3.16 ;
        RECT 1.36 2.235 2.06 2.435 ;
        RECT 1.36 0.605 1.625 1.31 ;
        RECT 1.36 0.605 1.53 2.435 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.89 2.555 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.91 -0.22 2.17 1.31 ;
        RECT 0.89 -0.22 1.15 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.25 2.08 0.51 2.88 ;
      RECT 0.25 2.08 1.15 2.26 ;
      RECT 0.89 1.05 1.15 2.26 ;
      RECT 0.25 1.05 1.15 1.31 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2b_1

MACRO sg13g2_nor2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2b_2 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 1.54 3 1.915 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.4 0.63 0.98 ;
    END
  END B_N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9728 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 1.16 2.6 1.36 ;
        RECT 2.34 0.72 2.6 1.36 ;
        RECT 1.83 2.08 2.09 2.68 ;
        RECT 1.36 2.08 2.09 2.285 ;
        RECT 1.36 0.72 1.58 2.285 ;
        RECT 1.32 0.72 1.58 1.42 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.85 2.22 3.11 4 ;
        RECT 0.81 2.22 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.85 -0.22 3.11 1.34 ;
        RECT 1.83 -0.22 2.09 0.98 ;
        RECT 0.81 -0.22 1.07 1.34 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.32 2.92 2.6 3.16 ;
      RECT 2.34 2.22 2.6 3.16 ;
      RECT 1.32 2.56 1.58 3.16 ;
      RECT 0.27 1.16 0.53 3.04 ;
      RECT 0.27 1.655 1.18 1.915 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2b_2

MACRO sg13g2_nor3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor3_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 1.515 0.62 1.85 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 1.515 1.58 1.85 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 1.515 2.06 1.85 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9814 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.965 2.22 2.225 3.13 ;
        RECT 0.945 1.06 2.225 1.22 ;
        RECT 1.965 0.62 2.225 1.22 ;
        RECT 0.945 2.38 2.225 2.665 ;
        RECT 0.945 0.62 1.205 1.22 ;
        RECT 0.945 0.62 1.12 2.665 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.375 2.205 0.635 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.455 -0.22 1.715 0.88 ;
        RECT 0.375 -0.22 0.635 1.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor3_1

MACRO sg13g2_nor3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor3_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 1.56 1.21 1.8 ;
        RECT 0.765 1.56 1.025 1.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.595 1.56 2.075 1.8 ;
        RECT 1.795 1.56 2.055 1.88 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.2 1.56 3.76 1.8 ;
        RECT 3.26 1.56 3.52 1.88 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2692 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.31 2.135 3.57 2.765 ;
        RECT 2.82 1.16 3.57 1.35 ;
        RECT 3.31 0.72 3.57 1.35 ;
        RECT 2.82 2.135 3.57 2.335 ;
        RECT 2.82 1.16 3.02 2.335 ;
        RECT 2.29 1.56 3.02 1.8 ;
        RECT 2.29 0.72 2.55 1.8 ;
        RECT 0.76 1.16 2.55 1.34 ;
        RECT 0.76 0.72 1.02 1.34 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 1.27 2.56 1.53 4 ;
        RECT 0.25 2.22 0.51 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.325 0.22 ;
        RECT 3.82 -0.22 4.08 1.32 ;
        RECT 2.8 -0.22 3.06 0.98 ;
        RECT 1.27 -0.22 2.04 0.98 ;
        RECT 0.25 -0.22 0.51 1.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.78 2.945 4.08 3.16 ;
      RECT 3.82 2.165 4.08 3.16 ;
      RECT 2.8 2.56 3.06 3.16 ;
      RECT 1.78 2.56 2.04 3.16 ;
      RECT 0.76 2.165 1.02 3.16 ;
      RECT 2.29 2.165 2.55 2.765 ;
      RECT 0.76 2.165 2.55 2.38 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor3_2

MACRO sg13g2_nor4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor4_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 1.455 0.63 1.905 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 1.455 1.23 1.735 ;
        RECT 0.835 1.455 1.08 1.905 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.41 1.455 1.72 1.735 ;
        RECT 1.3 1.905 1.58 2.335 ;
        RECT 1.41 1.455 1.58 2.335 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 1.455 2.32 1.905 ;
        RECT 1.8 2.335 2.06 2.74 ;
        RECT 1.9 1.455 2.06 2.74 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.28 2.22 2.7 3.16 ;
        RECT 2.505 1.05 2.7 3.16 ;
        RECT 0.81 1.05 2.7 1.21 ;
        RECT 1.83 0.61 2.09 1.21 ;
        RECT 0.81 0.61 1.07 1.21 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 0.3 2.22 0.56 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.34 -0.22 2.6 0.87 ;
        RECT 1.32 -0.22 1.58 0.87 ;
        RECT 0.3 -0.22 0.56 1.21 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor4_1

MACRO sg13g2_nor4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor4_2 0 0 ;
  SIZE 5.76 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.59 1.56 1.19 1.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.56 2.72 1.88 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.14 1.56 3.74 1.88 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5504 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.84 1.52 5.485 1.84 ;
        RECT 4.84 0.72 5.1 2.82 ;
        RECT 0.76 1.16 5.1 1.35 ;
        RECT 3.31 0.72 3.57 1.35 ;
        RECT 2.29 0.72 2.55 1.35 ;
        RECT 0.76 0.72 1.02 1.35 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 5.76 0.22 ;
        RECT 5.35 -0.22 5.61 1.32 ;
        RECT 3.82 -0.22 4.59 0.98 ;
        RECT 2.8 -0.22 3.06 0.98 ;
        RECT 1.27 -0.22 2.04 0.98 ;
        RECT 0.25 -0.22 0.51 1.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 5.76 4 ;
        RECT 1.27 2.56 1.53 4 ;
        RECT 0.25 2.22 0.51 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.025 1.56 4.64 1.88 ;
    END
  END D
  OBS
    LAYER Metal1 ;
      RECT 4.33 3 5.61 3.16 ;
      RECT 5.35 2.08 5.61 3.16 ;
      RECT 4.33 2.18 4.59 3.16 ;
      RECT 3.31 2.18 3.57 2.82 ;
      RECT 3.31 2.18 4.59 2.38 ;
      RECT 1.78 3 4.08 3.18 ;
      RECT 3.82 2.56 4.08 3.18 ;
      RECT 2.8 2.22 3.06 3.18 ;
      RECT 1.78 2.56 2.04 3.18 ;
      RECT 0.76 2.18 1.02 3.16 ;
      RECT 2.29 2.18 2.55 2.82 ;
      RECT 0.76 2.18 2.55 2.38 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor4_2

MACRO sg13g2_o21ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_o21ai_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 1.75 1.635 2.01 ;
        RECT 1.32 1.43 1.56 2.01 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.72 2.66 1.98 4 ;
        RECT 0.13 2.32 0.39 4 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.19 2.27 2.09 2.48 ;
        RECT 1.87 0.57 2.09 2.48 ;
        RECT 1.72 0.57 2.09 1.22 ;
        RECT 1.19 2.27 1.45 3.26 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.66 -0.22 0.92 0.84 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.24 1.43 0.6 2.01 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 1.43 1.08 2.01 ;
    END
  END A2
  OBS
    LAYER Metal1 ;
      RECT 0.13 1.06 1.45 1.245 ;
      RECT 1.19 0.57 1.45 1.245 ;
      RECT 0.13 0.57 0.39 1.245 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_o21ai_1

MACRO sg13g2_or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or2_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.315 -0.22 1.575 0.76 ;
        RECT 0.26 -0.22 0.52 0.76 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.3 2.34 1.56 4 ;
    END
  END VDD
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6492 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 2.34 2.15 3.28 ;
        RECT 1.955 0.5 2.15 3.28 ;
        RECT 1.825 0.5 2.15 1.1 ;
    END
  END X
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 2.13 1.08 2.65 ;
        RECT 0.625 2.13 1.08 2.37 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.635 1.255 1.895 ;
        RECT 0.84 1.495 1.08 1.895 ;
    END
  END A
  OBS
    LAYER Metal1 ;
      RECT 0.26 2.68 0.52 3.28 ;
      RECT 0.26 0.94 0.445 3.28 ;
      RECT 1.445 1.315 1.77 1.58 ;
      RECT 1.445 0.94 1.635 1.58 ;
      RECT 0.26 0.94 1.635 1.12 ;
      RECT 0.77 0.5 1.03 1.12 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or2_1

MACRO sg13g2_or2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.405 -0.22 2.665 1.1 ;
        RECT 1.275 -0.22 1.535 0.76 ;
        RECT 0.22 -0.22 0.48 0.76 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.405 2.34 2.665 4 ;
        RECT 1.27 2.34 1.53 4 ;
    END
  END VDD
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.837 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 2.34 2.05 3.28 ;
        RECT 1.885 0.5 2.05 3.28 ;
        RECT 1.785 0.5 2.05 1.1 ;
    END
  END X
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 2.13 1.085 2.88 ;
        RECT 0.585 2.13 1.085 2.35 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.635 1.215 1.895 ;
        RECT 0.84 1.335 1.085 1.895 ;
    END
  END A
  OBS
    LAYER Metal1 ;
      RECT 0.22 2.53 0.48 3.28 ;
      RECT 0.22 0.945 0.405 3.28 ;
      RECT 1.425 1.315 1.705 1.58 ;
      RECT 1.425 0.945 1.595 1.58 ;
      RECT 0.22 0.945 1.595 1.125 ;
      RECT 0.73 0.5 0.99 1.125 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or2_2

MACRO sg13g2_or3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or3_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.74 1.505 2.07 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.505 1.56 1.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.505 0.835 1.9 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.22 3.05 3.16 ;
        RECT 2.89 0.605 3.05 3.16 ;
        RECT 2.76 0.605 3.05 1.215 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 1.85 2.475 2.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.255 -0.22 2.515 0.87 ;
        RECT 0.895 -0.22 1.155 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.385 2.09 0.645 3.04 ;
      RECT 0.385 2.09 2.515 2.295 ;
      RECT 2.345 1.115 2.515 2.295 ;
      RECT 2.345 1.52 2.71 1.85 ;
      RECT 0.385 1.115 2.515 1.325 ;
      RECT 0.385 1.11 1.965 1.325 ;
      RECT 1.445 0.61 1.965 1.325 ;
      RECT 0.385 0.61 0.645 1.325 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or3_1

MACRO sg13g2_or3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or3_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.74 1.505 2.07 1.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.505 1.56 1.935 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.505 0.835 1.935 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7142 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.89 1.485 3.64 1.855 ;
        RECT 2.7 2.215 3.05 3.16 ;
        RECT 2.89 0.605 3.05 3.16 ;
        RECT 2.76 0.605 3.05 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.27 2.22 3.53 4 ;
        RECT 1.85 2.475 2.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.285 -0.22 3.545 1.21 ;
        RECT 2.255 -0.22 2.515 0.87 ;
        RECT 0.895 -0.22 1.155 0.89 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.385 2.12 0.645 3.04 ;
      RECT 0.385 2.12 2.515 2.295 ;
      RECT 2.345 1.115 2.515 2.295 ;
      RECT 2.345 1.57 2.71 1.85 ;
      RECT 0.385 1.115 2.515 1.325 ;
      RECT 0.385 1.11 1.965 1.325 ;
      RECT 1.445 0.61 1.965 1.325 ;
      RECT 0.385 0.61 0.645 1.325 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or3_2

MACRO sg13g2_or4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or4_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.545 2.605 1.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 1.545 2.045 1.935 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 1.545 1.56 1.935 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.32 1.545 0.875 1.935 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 2.095 3.5 3.145 ;
        RECT 3.34 0.62 3.5 3.145 ;
        RECT 3.18 0.62 3.5 1.295 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.645 2.585 2.905 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.635 -0.22 2.895 1.01 ;
        RECT 1.455 -0.22 1.715 1 ;
        RECT 0.38 -0.22 0.64 1.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.38 2.555 0.64 3.16 ;
      RECT 0.38 2.555 2.36 2.75 ;
      RECT 2.2 2.19 2.36 2.75 ;
      RECT 2.2 2.19 2.955 2.38 ;
      RECT 2.785 1.195 2.955 2.38 ;
      RECT 2.785 1.52 3.16 1.85 ;
      RECT 2.785 1.195 2.995 1.85 ;
      RECT 0.89 1.195 2.995 1.365 ;
      RECT 2.115 0.855 2.375 1.365 ;
      RECT 0.89 0.855 1.15 1.365 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or4_1

MACRO sg13g2_or4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or4_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.545 2.605 1.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 1.545 2.045 1.97 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.18 1.545 1.57 1.97 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 1.545 0.875 1.935 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7681 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 2.22 3.5 3.16 ;
        RECT 3.34 0.61 3.5 3.16 ;
        RECT 3.18 0.61 3.5 1.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.72 2.22 3.98 4 ;
        RECT 2.645 2.585 2.905 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.69 -0.22 3.95 1.21 ;
        RECT 2.625 -0.22 2.885 1.01 ;
        RECT 1.455 -0.22 1.715 1.015 ;
        RECT 0.38 -0.22 0.64 1.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.38 2.19 0.64 3.16 ;
      RECT 0.38 2.19 2.955 2.38 ;
      RECT 2.785 1.195 2.955 2.38 ;
      RECT 2.785 1.52 3.16 1.85 ;
      RECT 2.785 1.195 2.995 1.85 ;
      RECT 0.89 1.195 2.995 1.365 ;
      RECT 2.115 0.8 2.375 1.365 ;
      RECT 0.89 0.8 1.15 1.365 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or4_2

MACRO sg13g2_sdfbbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfbbp_1 0 0 ;
  SIZE 16.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.145 0.59 16.535 3.12 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.59 2.005 14.95 3.135 ;
        RECT 14.78 0.61 14.95 3.135 ;
        RECT 14.52 0.61 14.95 1.19 ;
    END
  END Q_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.74 1.38 14.035 1.79 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.51 1.72 11.84 2 ;
        RECT 11.51 1.72 11.81 2.35 ;
        RECT 10.58 1.89 11.81 2.05 ;
        RECT 9.31 3.105 10.74 3.275 ;
        RECT 10.58 1.89 10.74 3.275 ;
        RECT 10.565 2.215 10.74 3.275 ;
        RECT 9.31 2.345 9.48 3.275 ;
        RECT 8.39 2.345 9.48 2.51 ;
        RECT 7.55 3.105 8.56 3.275 ;
        RECT 8.39 2.345 8.56 3.275 ;
        RECT 7.525 1.635 7.815 1.855 ;
        RECT 7.55 1.635 7.72 3.275 ;
    END
  END SET_B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal2 ;
      ANTENNAMAXAREACAR 1.167997 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.261974 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.68 1.62 2.05 2.055 ;
      LAYER Metal2 ;
        RECT 1.645 1.58 2.205 1.86 ;
      LAYER Via1 ;
        RECT 1.79 1.645 1.98 1.835 ;
    END
  END D
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2756 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 1.75 1.435 2.295 ;
    END
  END SCE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.51 1.355 0.84 2.325 ;
    END
  END SCD
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.885 1.38 4.34 1.85 ;
        RECT 3.92 1.155 4.34 1.85 ;
    END
  END CLK
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 16.8 4 ;
        RECT 15.645 2.455 15.905 4 ;
        RECT 14.055 2.885 14.315 4 ;
        RECT 12.765 2.88 13.025 4 ;
        RECT 10.925 3.055 11.57 4 ;
        RECT 8.815 2.695 9.075 4 ;
        RECT 6.915 2.34 7.175 4 ;
        RECT 4.46 2.56 4.72 4 ;
        RECT 2.92 2.88 3.18 4 ;
        RECT 0.85 2.88 1.11 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 16.8 0.22 ;
        RECT 15.675 -0.22 15.935 1.155 ;
        RECT 14.035 -0.22 14.295 1.14 ;
        RECT 11.34 -0.22 11.6 1.16 ;
        RECT 9.415 -0.22 9.59 1.175 ;
        RECT 7.01 -0.22 7.27 0.745 ;
        RECT 4.26 -0.22 4.46 0.635 ;
        RECT 2.185 -0.22 2.445 1.095 ;
        RECT 0.34 -0.22 0.6 1.055 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 15.17 1.555 15.375 3.07 ;
      RECT 15.17 1.555 15.645 1.885 ;
      RECT 15.17 0.705 15.355 3.07 ;
      RECT 11.93 2.66 12.205 3.145 ;
      RECT 11.99 2.195 12.205 3.145 ;
      RECT 10.92 2.66 12.205 2.87 ;
      RECT 10.92 2.23 11.25 2.87 ;
      RECT 11.99 2.485 14.375 2.645 ;
      RECT 14.215 1.42 14.375 2.645 ;
      RECT 11.99 2.195 12.67 2.645 ;
      RECT 12.51 0.875 12.67 2.645 ;
      RECT 14.215 1.42 14.55 1.75 ;
      RECT 12.34 0.875 12.67 1.125 ;
      RECT 13.34 1.975 13.795 2.305 ;
      RECT 13.34 0.93 13.5 2.305 ;
      RECT 12.9 1.38 13.5 1.865 ;
      RECT 13.34 0.93 13.815 1.14 ;
      RECT 12.87 0.515 13.13 1.17 ;
      RECT 11.85 0.515 12.11 1.155 ;
      RECT 11.85 0.515 13.13 0.695 ;
      RECT 9.83 2.31 10.38 2.895 ;
      RECT 10.21 0.935 10.38 2.895 ;
      RECT 12.05 1.345 12.33 1.75 ;
      RECT 10.21 1.55 11.25 1.71 ;
      RECT 11.085 1.345 11.25 1.71 ;
      RECT 10.21 0.935 10.44 1.71 ;
      RECT 11.085 1.345 12.33 1.525 ;
      RECT 9.71 1.755 10.03 2.125 ;
      RECT 9.71 1.535 9.93 2.125 ;
      RECT 9.77 0.455 9.93 2.125 ;
      RECT 10.645 0.455 10.905 1.36 ;
      RECT 9.77 0.455 10.905 0.615 ;
      RECT 7.925 2 8.16 2.905 ;
      RECT 7.925 2 9.47 2.16 ;
      RECT 9.075 1.535 9.47 2.16 ;
      RECT 6.77 0.955 6.975 1.65 ;
      RECT 9.075 0.955 9.235 2.16 ;
      RECT 6.77 0.955 9.235 1.115 ;
      RECT 8.255 0.87 8.515 1.115 ;
      RECT 8.795 0.52 9.055 0.775 ;
      RECT 7.71 0.52 8.005 0.775 ;
      RECT 7.71 0.52 9.055 0.68 ;
      RECT 6.065 2.465 6.58 2.67 ;
      RECT 6.42 0.825 6.58 2.67 ;
      RECT 6.42 1.995 7.33 2.16 ;
      RECT 7.16 1.295 7.33 2.16 ;
      RECT 8.04 1.295 8.37 1.785 ;
      RECT 7.16 1.295 8.37 1.455 ;
      RECT 5.955 0.825 6.58 0.985 ;
      RECT 5.955 0.725 6.22 0.985 ;
      RECT 5.585 2.075 5.785 2.92 ;
      RECT 1.88 2.255 2.14 2.845 ;
      RECT 1.88 2.255 2.495 2.455 ;
      RECT 2.29 1.28 2.495 2.455 ;
      RECT 5.585 2.075 6.24 2.235 ;
      RECT 6.08 1.225 6.24 2.235 ;
      RECT 1.36 1.28 2.85 1.44 ;
      RECT 2.67 0.455 2.85 1.44 ;
      RECT 5.54 1.225 6.24 1.385 ;
      RECT 1.36 0.875 1.62 1.44 ;
      RECT 5.54 0.7 5.73 1.385 ;
      RECT 3.92 0.815 5.73 0.975 ;
      RECT 5.425 0.7 5.73 0.975 ;
      RECT 3.92 0.455 4.08 0.975 ;
      RECT 2.67 0.455 4.08 0.625 ;
      RECT 4.985 2.22 5.245 3.16 ;
      RECT 5.19 1.155 5.36 2.49 ;
      RECT 5.19 1.58 5.9 1.88 ;
      RECT 4.77 1.155 5.36 1.335 ;
      RECT 3.95 2.04 4.21 3.16 ;
      RECT 3.535 2.04 4.7 2.21 ;
      RECT 4.53 1.54 4.7 2.21 ;
      RECT 3.535 0.87 3.695 2.21 ;
      RECT 4.53 1.54 5.005 1.87 ;
      RECT 3.535 0.87 3.74 1.21 ;
      RECT 3.43 2.47 3.69 3.14 ;
      RECT 3.03 2.47 3.69 2.64 ;
      RECT 3.03 0.885 3.215 2.64 ;
      RECT 2.675 2.065 3.215 2.325 ;
      RECT 1.355 3.105 2.66 3.275 ;
      RECT 2.4 2.88 2.66 3.275 ;
      RECT 0.34 2.505 0.6 3.14 ;
      RECT 1.355 2.505 1.555 3.275 ;
      RECT 0.34 2.505 1.555 2.675 ;
      RECT 8.58 1.38 8.885 1.785 ;
    LAYER Via1 ;
      RECT 13.09 1.595 13.28 1.785 ;
      RECT 8.685 1.52 8.875 1.71 ;
    LAYER Metal2 ;
      RECT 8.635 1.455 9 1.9 ;
      RECT 13.03 1.47 13.32 1.865 ;
      RECT 8.635 1.58 13.32 1.78 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfbbp_1

MACRO sg13g2_sdfrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfrbp_1 0 0 ;
  SIZE 18.24 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7 1.51 7.55 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 18.24 0.22 ;
        RECT 17.3 -0.22 17.555 1.21 ;
        RECT 16.27 -0.22 16.53 0.85 ;
        RECT 14.36 -0.22 14.62 0.885 ;
        RECT 7.035 -0.22 7.295 0.915 ;
        RECT 5.94 -0.22 6.2 0.885 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 18.24 4 ;
        RECT 17.3 2.235 17.56 4 ;
        RECT 16.27 1.98 16.53 4 ;
        RECT 15.25 2.46 15.51 4 ;
        RECT 7.745 2.86 7.915 4 ;
        RECT 5.015 2.215 5.27 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.92 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END SCD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 17.81 0.595 18.07 3.175 ;
        RECT 17.525 1.51 18.07 1.855 ;
        RECT 17.805 0.595 18.07 1.855 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.165 1.335 11.79 1.935 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.4 2.535 1.92 ;
    END
  END D
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6842 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.76 1.06 16.52 1.45 ;
        RECT 15.76 0.59 16.02 3.06 ;
    END
  END Q_N
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.5 1.105 1.87 ;
    END
  END SCE
  OBS
    LAYER Metal1 ;
      RECT 16.78 0.59 17.04 2.92 ;
      RECT 16.775 0.59 17.04 1.98 ;
      RECT 16.775 1.535 17.2 1.795 ;
      RECT 14.71 2.1 14.97 2.495 ;
      RECT 13.93 2.1 15.53 2.26 ;
      RECT 15.37 0.625 15.53 2.26 ;
      RECT 13.93 1.655 14.185 2.26 ;
      RECT 15.18 0.625 15.53 0.885 ;
      RECT 13.255 2.125 13.46 2.5 ;
      RECT 13.255 2.125 13.75 2.295 ;
      RECT 13.59 1.145 13.75 2.295 ;
      RECT 14.965 1.275 15.19 1.665 ;
      RECT 13.59 1.275 15.19 1.465 ;
      RECT 12.76 1.145 13.77 1.315 ;
      RECT 14.71 3.025 14.98 3.285 ;
      RECT 9.655 3.025 9.915 3.285 ;
      RECT 9.655 3.075 14.98 3.235 ;
      RECT 12.31 0.805 12.48 1.31 ;
      RECT 12.31 0.805 14.11 0.965 ;
      RECT 13.85 0.625 14.11 0.965 ;
      RECT 6 2.64 6.74 2.9 ;
      RECT 6 1.17 6.16 2.9 ;
      RECT 12.545 1.555 12.735 2.45 ;
      RECT 7.735 1.755 8.015 1.965 ;
      RECT 7.735 1.17 7.895 1.965 ;
      RECT 11.97 1.555 12.735 1.725 ;
      RECT 11.97 0.44 12.13 1.725 ;
      RECT 6 1.17 7.895 1.33 ;
      RECT 7.505 0.44 7.675 1.33 ;
      RECT 6.52 0.815 6.78 1.33 ;
      RECT 13.34 0.44 13.6 0.625 ;
      RECT 7.505 0.44 13.6 0.605 ;
      RECT 10.225 2.63 13.075 2.79 ;
      RECT 12.915 1.51 13.075 2.79 ;
      RECT 10.225 2.06 10.585 2.79 ;
      RECT 9.82 2.15 10.585 2.41 ;
      RECT 9.955 2.06 10.585 2.41 ;
      RECT 9.955 1.135 10.215 2.41 ;
      RECT 12.915 1.51 13.4 1.77 ;
      RECT 10.765 2.145 12.325 2.37 ;
      RECT 12.065 2.075 12.325 2.37 ;
      RECT 10.765 0.855 10.925 2.37 ;
      RECT 10.45 1.54 10.925 1.87 ;
      RECT 11.555 0.81 11.79 1.07 ;
      RECT 10.765 0.855 11.79 1.025 ;
      RECT 9.43 1.44 9.695 1.7 ;
      RECT 9.485 1.3 9.695 1.7 ;
      RECT 9.485 0.785 9.665 1.7 ;
      RECT 7.965 0.785 9.665 0.96 ;
      RECT 5.59 3.08 7.565 3.24 ;
      RECT 7.405 2.52 7.565 3.24 ;
      RECT 8.255 2.985 9.425 3.145 ;
      RECT 9.09 2.685 9.425 3.145 ;
      RECT 5.59 2.24 5.78 3.24 ;
      RECT 8.255 2.52 8.415 3.145 ;
      RECT 9.09 1.17 9.25 3.145 ;
      RECT 7.405 2.52 8.415 2.68 ;
      RECT 5.52 2.24 5.78 2.52 ;
      RECT 5.59 0.645 5.75 3.24 ;
      RECT 8.185 1.225 8.445 1.64 ;
      RECT 8.265 1.17 9.25 1.33 ;
      RECT 5.01 0.645 5.75 0.84 ;
      RECT 7.045 2.145 7.225 2.9 ;
      RECT 8.69 1.51 8.875 2.805 ;
      RECT 7.045 2.145 8.875 2.315 ;
      RECT 6.385 2.145 8.875 2.305 ;
      RECT 6.385 1.705 6.645 2.305 ;
      RECT 8.69 1.51 8.91 1.81 ;
      RECT 4.135 2.04 4.59 3.2 ;
      RECT 4.4 0.57 4.59 3.2 ;
      RECT 5.055 1.445 5.315 1.75 ;
      RECT 4.4 1.445 5.315 1.7 ;
      RECT 4.315 0.57 4.59 1.21 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.855 2.345 2.56 2.505 ;
      RECT 1.855 2.08 2.015 2.505 ;
      RECT 1.285 2.08 2.015 2.26 ;
      RECT 1.285 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.22 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.285 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.295 2.28 0.575 2.88 ;
      RECT 0.295 2.44 1.64 2.6 ;
      RECT 0.295 0.8 0.455 2.88 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.295 0.8 0.575 1.06 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfrbp_1

MACRO sg13g2_sdfrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfrbp_2 0 0 ;
  SIZE 19.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7 1.51 7.55 1.965 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 19.2 0.22 ;
        RECT 18.735 -0.22 19.01 0.84 ;
        RECT 17.73 -0.22 17.99 1.21 ;
        RECT 16.71 -0.22 16.97 0.85 ;
        RECT 15.71 -0.22 15.95 0.85 ;
        RECT 14.36 -0.22 14.62 0.885 ;
        RECT 7.035 -0.22 7.295 0.915 ;
        RECT 5.94 -0.22 6.2 0.885 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 19.2 4 ;
        RECT 18.38 2.085 18.64 4 ;
        RECT 17.355 2.085 17.615 4 ;
        RECT 16.27 1.98 16.53 4 ;
        RECT 15.25 2.46 15.51 4 ;
        RECT 7.745 2.86 7.915 4 ;
        RECT 5.015 2.215 5.27 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.92 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END SCD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7124 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 18.24 1.045 19.01 1.49 ;
        RECT 17.99 1.515 18.5 1.775 ;
        RECT 18.24 0.595 18.5 1.775 ;
        RECT 17.865 2.085 18.16 3.175 ;
        RECT 17.99 1.515 18.16 3.175 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.165 1.335 11.79 1.935 ;
    END
  END CLK
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.5 1.105 1.87 ;
    END
  END SCE
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.76 1.52 16.52 1.74 ;
        RECT 16.14 0.99 16.52 1.74 ;
        RECT 16.195 0.59 16.46 1.74 ;
        RECT 15.76 1.52 16.02 3.06 ;
    END
  END Q_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.4 2.535 1.92 ;
    END
  END D
  OBS
    LAYER Metal1 ;
      RECT 16.78 1.98 17.16 2.92 ;
      RECT 16.99 1.535 17.16 2.92 ;
      RECT 16.99 1.535 17.785 1.795 ;
      RECT 17.2 0.59 17.485 1.795 ;
      RECT 14.71 2.1 14.97 2.495 ;
      RECT 13.93 2.1 15.53 2.26 ;
      RECT 15.37 0.625 15.53 2.26 ;
      RECT 13.93 1.655 14.185 2.26 ;
      RECT 15.18 0.625 15.53 0.885 ;
      RECT 13.255 2.125 13.46 2.5 ;
      RECT 13.255 2.125 13.75 2.295 ;
      RECT 13.59 1.145 13.75 2.295 ;
      RECT 14.965 1.275 15.19 1.665 ;
      RECT 13.59 1.275 15.19 1.465 ;
      RECT 12.76 1.145 13.77 1.315 ;
      RECT 14.71 3.025 14.98 3.285 ;
      RECT 9.655 3.025 9.915 3.285 ;
      RECT 9.655 3.075 14.98 3.235 ;
      RECT 12.31 0.805 12.48 1.31 ;
      RECT 12.31 0.805 14.11 0.965 ;
      RECT 13.85 0.625 14.11 0.965 ;
      RECT 6 2.64 6.74 2.9 ;
      RECT 6 1.17 6.16 2.9 ;
      RECT 12.545 1.555 12.735 2.45 ;
      RECT 7.735 1.755 8.015 1.965 ;
      RECT 7.735 1.17 7.895 1.965 ;
      RECT 11.97 1.555 12.735 1.725 ;
      RECT 11.97 0.44 12.13 1.725 ;
      RECT 6 1.17 7.895 1.33 ;
      RECT 7.505 0.44 7.675 1.33 ;
      RECT 6.52 0.815 6.78 1.33 ;
      RECT 13.34 0.44 13.6 0.625 ;
      RECT 7.505 0.44 13.6 0.605 ;
      RECT 10.225 2.63 13.075 2.79 ;
      RECT 12.915 1.51 13.075 2.79 ;
      RECT 10.225 2.06 10.585 2.79 ;
      RECT 9.82 2.15 10.585 2.41 ;
      RECT 9.955 2.06 10.585 2.41 ;
      RECT 9.955 1.135 10.215 2.41 ;
      RECT 12.915 1.51 13.4 1.77 ;
      RECT 10.765 2.145 12.325 2.37 ;
      RECT 12.065 2.075 12.325 2.37 ;
      RECT 10.765 0.855 10.925 2.37 ;
      RECT 10.45 1.54 10.925 1.87 ;
      RECT 11.555 0.81 11.79 1.07 ;
      RECT 10.765 0.855 11.79 1.025 ;
      RECT 9.43 1.44 9.695 1.7 ;
      RECT 9.485 1.3 9.695 1.7 ;
      RECT 9.485 0.785 9.665 1.7 ;
      RECT 7.965 0.785 9.665 0.96 ;
      RECT 5.59 3.08 7.565 3.24 ;
      RECT 7.405 2.52 7.565 3.24 ;
      RECT 8.255 2.985 9.425 3.145 ;
      RECT 9.09 2.685 9.425 3.145 ;
      RECT 5.59 2.24 5.78 3.24 ;
      RECT 8.255 2.52 8.415 3.145 ;
      RECT 9.09 1.17 9.25 3.145 ;
      RECT 7.405 2.52 8.415 2.68 ;
      RECT 5.52 2.24 5.78 2.52 ;
      RECT 5.59 0.645 5.75 3.24 ;
      RECT 8.185 1.225 8.445 1.64 ;
      RECT 8.265 1.17 9.25 1.33 ;
      RECT 5.01 0.645 5.75 0.84 ;
      RECT 7.045 2.145 7.225 2.9 ;
      RECT 8.69 1.51 8.875 2.805 ;
      RECT 7.045 2.145 8.875 2.315 ;
      RECT 6.385 2.145 8.875 2.305 ;
      RECT 6.385 1.705 6.645 2.305 ;
      RECT 8.69 1.51 8.91 1.81 ;
      RECT 4.135 2.04 4.59 3.2 ;
      RECT 4.4 0.57 4.59 3.2 ;
      RECT 4.4 1.49 5.315 1.75 ;
      RECT 4.315 0.57 4.59 1.21 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.855 2.345 2.56 2.505 ;
      RECT 1.855 2.08 2.015 2.505 ;
      RECT 1.285 2.08 2.015 2.26 ;
      RECT 1.285 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.22 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.285 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.295 2.28 0.575 2.88 ;
      RECT 0.295 2.44 1.64 2.6 ;
      RECT 0.295 0.8 0.455 2.88 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.295 0.8 0.575 1.06 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfrbp_2

MACRO sg13g2_sdfrbpq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfrbpq_1 0 0 ;
  SIZE 16.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.055 1 16.57 1.465 ;
        RECT 16.28 0.59 16.54 3.02 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.165 1.335 11.79 1.935 ;
    END
  END CLK
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7 1.51 7.55 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.92 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END SCD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.4 2.535 1.92 ;
    END
  END D
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.5 1.105 1.87 ;
    END
  END SCE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 16.8 0.22 ;
        RECT 15.77 -0.22 16.03 0.81 ;
        RECT 14.36 -0.22 14.62 0.885 ;
        RECT 7.035 -0.22 7.295 0.915 ;
        RECT 5.94 -0.22 6.2 0.885 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 16.8 4 ;
        RECT 15.77 2.08 16.03 4 ;
        RECT 15.25 2.46 15.51 4 ;
        RECT 7.745 2.86 7.915 4 ;
        RECT 5.015 2.215 5.27 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      RECT 14.71 2.1 14.97 2.495 ;
      RECT 13.93 2.1 15.53 2.26 ;
      RECT 15.37 0.625 15.53 2.26 ;
      RECT 13.93 1.655 14.185 2.26 ;
      RECT 15.37 1.61 15.9 1.84 ;
      RECT 15.18 0.625 15.53 0.885 ;
      RECT 13.255 2.125 13.46 2.5 ;
      RECT 13.255 2.125 13.75 2.295 ;
      RECT 13.59 1.145 13.75 2.295 ;
      RECT 14.965 1.275 15.19 1.665 ;
      RECT 13.59 1.275 15.19 1.465 ;
      RECT 12.76 1.145 13.77 1.315 ;
      RECT 14.71 3.025 14.98 3.285 ;
      RECT 9.655 3.025 9.915 3.285 ;
      RECT 9.655 3.075 14.98 3.235 ;
      RECT 12.31 0.805 12.48 1.31 ;
      RECT 12.31 0.805 14.11 0.965 ;
      RECT 13.85 0.625 14.11 0.965 ;
      RECT 6 2.64 6.74 2.9 ;
      RECT 6 1.17 6.16 2.9 ;
      RECT 12.545 1.555 12.735 2.45 ;
      RECT 7.735 1.755 8.015 1.965 ;
      RECT 7.735 1.17 7.895 1.965 ;
      RECT 11.97 1.555 12.735 1.725 ;
      RECT 11.97 0.44 12.13 1.725 ;
      RECT 6 1.17 7.895 1.33 ;
      RECT 7.505 0.44 7.675 1.33 ;
      RECT 6.52 0.815 6.78 1.33 ;
      RECT 13.34 0.44 13.6 0.625 ;
      RECT 7.505 0.44 13.6 0.605 ;
      RECT 10.225 2.63 13.075 2.79 ;
      RECT 12.915 1.51 13.075 2.79 ;
      RECT 10.225 2.06 10.585 2.79 ;
      RECT 9.82 2.15 10.585 2.41 ;
      RECT 9.955 2.06 10.585 2.41 ;
      RECT 9.955 1.135 10.215 2.41 ;
      RECT 12.915 1.51 13.4 1.77 ;
      RECT 10.765 2.145 12.325 2.37 ;
      RECT 12.065 2.075 12.325 2.37 ;
      RECT 10.765 0.855 10.925 2.37 ;
      RECT 10.45 1.54 10.925 1.87 ;
      RECT 11.555 0.81 11.79 1.07 ;
      RECT 10.765 0.855 11.79 1.025 ;
      RECT 9.43 1.44 9.695 1.7 ;
      RECT 9.485 1.3 9.695 1.7 ;
      RECT 9.485 0.785 9.665 1.7 ;
      RECT 7.965 0.785 9.665 0.96 ;
      RECT 5.59 3.08 7.565 3.24 ;
      RECT 7.405 2.52 7.565 3.24 ;
      RECT 8.255 2.985 9.425 3.145 ;
      RECT 9.09 2.685 9.425 3.145 ;
      RECT 5.59 2.24 5.78 3.24 ;
      RECT 8.255 2.52 8.415 3.145 ;
      RECT 9.09 1.17 9.25 3.145 ;
      RECT 7.405 2.52 8.415 2.68 ;
      RECT 5.52 2.24 5.78 2.52 ;
      RECT 5.59 0.645 5.75 3.24 ;
      RECT 8.185 1.225 8.445 1.64 ;
      RECT 8.265 1.17 9.25 1.33 ;
      RECT 5.01 0.645 5.75 0.84 ;
      RECT 7.045 2.145 7.225 2.9 ;
      RECT 8.69 1.51 8.875 2.805 ;
      RECT 7.045 2.145 8.875 2.315 ;
      RECT 6.385 2.145 8.875 2.305 ;
      RECT 6.385 1.705 6.645 2.305 ;
      RECT 8.69 1.51 8.91 1.81 ;
      RECT 4.135 2.04 4.59 3.2 ;
      RECT 4.4 0.57 4.59 3.2 ;
      RECT 5.055 1.445 5.315 1.75 ;
      RECT 4.4 1.445 5.315 1.7 ;
      RECT 4.315 0.57 4.59 1.21 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.855 2.345 2.56 2.505 ;
      RECT 1.855 2.08 2.015 2.505 ;
      RECT 1.285 2.08 2.015 2.26 ;
      RECT 1.285 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.22 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.285 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.295 2.28 0.575 2.88 ;
      RECT 0.295 2.44 1.64 2.6 ;
      RECT 0.295 0.8 0.455 2.88 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.295 0.8 0.575 1.06 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfrbpq_1

MACRO sg13g2_sdfrbpq_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfrbpq_2 0 0 ;
  SIZE 17.28 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.86 1.52 16.52 1.74 ;
        RECT 16.14 0.99 16.52 1.74 ;
        RECT 16.195 0.59 16.46 1.74 ;
        RECT 15.76 2.085 16.02 3.06 ;
        RECT 15.86 1.52 16.02 3.06 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.165 1.335 11.79 1.935 ;
    END
  END CLK
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.905 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.762515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7 1.51 7.55 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1.03 3.015 1.92 ;
        RECT 1.71 1.03 3.015 1.2 ;
        RECT 1.63 1.47 1.89 1.73 ;
        RECT 1.71 1.03 1.89 1.73 ;
    END
  END SCD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 1.4 2.535 1.92 ;
    END
  END D
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.5 1.105 1.87 ;
    END
  END SCE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 17.28 4 ;
        RECT 16.27 2.1 16.53 4 ;
        RECT 15.25 2.46 15.51 4 ;
        RECT 7.745 2.86 7.915 4 ;
        RECT 5.015 2.215 5.27 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.78 1.235 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 17.28 0.22 ;
        RECT 16.71 -0.22 16.97 1.195 ;
        RECT 15.71 -0.22 15.95 1.195 ;
        RECT 14.36 -0.22 14.62 0.885 ;
        RECT 7.035 -0.22 7.295 0.915 ;
        RECT 5.94 -0.22 6.2 0.885 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 14.71 2.1 14.97 2.495 ;
      RECT 13.93 2.1 15.53 2.26 ;
      RECT 15.37 0.625 15.53 2.26 ;
      RECT 13.93 1.655 14.185 2.26 ;
      RECT 15.37 1.575 15.68 1.835 ;
      RECT 15.18 0.625 15.53 0.885 ;
      RECT 13.255 2.125 13.46 2.5 ;
      RECT 13.255 2.125 13.75 2.295 ;
      RECT 13.59 1.145 13.75 2.295 ;
      RECT 14.915 1.275 15.175 1.665 ;
      RECT 13.59 1.275 15.175 1.465 ;
      RECT 12.76 1.145 13.77 1.315 ;
      RECT 14.71 3.025 14.98 3.285 ;
      RECT 9.655 3.025 9.915 3.285 ;
      RECT 9.655 3.075 14.98 3.235 ;
      RECT 12.31 0.805 12.48 1.31 ;
      RECT 12.31 0.805 14.11 0.965 ;
      RECT 13.85 0.625 14.11 0.965 ;
      RECT 6 2.64 6.74 2.9 ;
      RECT 6 1.17 6.16 2.9 ;
      RECT 12.545 1.555 12.735 2.45 ;
      RECT 7.735 1.755 8.015 1.965 ;
      RECT 7.735 1.17 7.895 1.965 ;
      RECT 11.97 1.555 12.735 1.725 ;
      RECT 11.97 0.44 12.13 1.725 ;
      RECT 6 1.17 7.895 1.33 ;
      RECT 7.505 0.44 7.675 1.33 ;
      RECT 6.52 0.815 6.78 1.33 ;
      RECT 13.34 0.44 13.6 0.625 ;
      RECT 7.505 0.44 13.6 0.605 ;
      RECT 10.225 2.63 13.075 2.79 ;
      RECT 12.915 1.51 13.075 2.79 ;
      RECT 10.225 2.06 10.585 2.79 ;
      RECT 9.82 2.15 10.585 2.41 ;
      RECT 9.955 2.06 10.585 2.41 ;
      RECT 9.955 1.135 10.215 2.41 ;
      RECT 12.915 1.51 13.4 1.77 ;
      RECT 10.765 2.145 12.325 2.37 ;
      RECT 12.065 2.075 12.325 2.37 ;
      RECT 10.765 0.855 10.925 2.37 ;
      RECT 10.45 1.54 10.925 1.87 ;
      RECT 11.555 0.81 11.79 1.07 ;
      RECT 10.765 0.855 11.79 1.025 ;
      RECT 9.43 1.44 9.695 1.7 ;
      RECT 9.485 1.3 9.695 1.7 ;
      RECT 9.485 0.785 9.665 1.7 ;
      RECT 7.965 0.785 9.665 0.96 ;
      RECT 5.59 3.08 7.565 3.24 ;
      RECT 7.405 2.52 7.565 3.24 ;
      RECT 8.255 2.985 9.425 3.145 ;
      RECT 9.09 2.685 9.425 3.145 ;
      RECT 5.59 2.24 5.78 3.24 ;
      RECT 8.255 2.52 8.415 3.145 ;
      RECT 9.09 1.17 9.25 3.145 ;
      RECT 7.405 2.52 8.415 2.68 ;
      RECT 5.52 2.24 5.78 2.52 ;
      RECT 5.59 0.645 5.75 3.24 ;
      RECT 8.185 1.225 8.445 1.64 ;
      RECT 8.265 1.17 9.25 1.33 ;
      RECT 5.01 0.645 5.75 0.84 ;
      RECT 7.045 2.145 7.225 2.9 ;
      RECT 8.69 1.51 8.875 2.805 ;
      RECT 7.045 2.145 8.875 2.315 ;
      RECT 6.385 2.145 8.875 2.305 ;
      RECT 6.385 1.705 6.645 2.305 ;
      RECT 8.69 1.51 8.91 1.81 ;
      RECT 4.135 2.04 4.59 3.2 ;
      RECT 4.4 0.57 4.59 3.2 ;
      RECT 4.4 1.49 5.315 1.75 ;
      RECT 4.315 0.57 4.59 1.21 ;
      RECT 2.3 2.345 2.56 2.945 ;
      RECT 1.855 2.345 2.56 2.505 ;
      RECT 1.855 2.08 2.015 2.505 ;
      RECT 1.285 2.08 2.015 2.26 ;
      RECT 1.285 0.61 1.45 2.26 ;
      RECT 3.945 1.52 4.22 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.285 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.44 1.64 3.295 ;
      RECT 0.295 2.28 0.575 2.88 ;
      RECT 0.295 2.44 1.64 2.6 ;
      RECT 0.295 0.8 0.455 2.88 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.295 0.8 0.575 1.06 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfrbpq_2

MACRO sg13g2_sighold
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sighold 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.57 3.17 1.925 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.555 -0.22 1.83 0.545 ;
    END
  END VSS
  PIN SH
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.204 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.955 2.045 2.41 ;
        RECT 0.585 1.765 2.045 2.025 ;
    END
  END SH
  OBS
    LAYER Metal1 ;
      RECT 0.175 1.325 0.405 2.41 ;
      RECT 0.175 1.325 1.245 1.585 ;
      RECT 0.175 0.955 0.395 2.41 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sighold

MACRO sg13g2_slgcp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_slgcp_1 0 0 ;
  SIZE 8.16 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.96 1.525 2.24 ;
        RECT 1.095 1.885 1.355 2.24 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 1.51 0.615 2.145 ;
    END
  END SCE
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3978 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.585 1.56 5.89 2 ;
    END
  END CLK
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.445 2.06 7.84 3.18 ;
        RECT 7.68 0.62 7.84 3.18 ;
        RECT 7.58 0.62 7.84 1.3 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.16 4 ;
        RECT 6.935 2.335 7.195 4 ;
        RECT 4.28 2.785 4.54 4 ;
        RECT 1.82 2.94 2.08 4 ;
        RECT 0.23 2.54 0.49 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.16 0.22 ;
        RECT 7.09 -0.22 7.275 1.22 ;
        RECT 5.66 -0.22 5.92 1.275 ;
        RECT 3.99 -0.22 4.15 0.91 ;
        RECT 1.28 -0.22 1.54 0.575 ;
        RECT 0.23 -0.22 0.49 1.165 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 6.455 1.94 6.65 3.075 ;
      RECT 6.455 1.94 6.9 2.11 ;
      RECT 6.74 0.71 6.9 2.11 ;
      RECT 6.74 1.52 7.5 1.85 ;
      RECT 6.74 0.71 6.91 1.85 ;
      RECT 6.485 0.71 6.91 1.27 ;
      RECT 4.79 2 5.05 3.065 ;
      RECT 4.79 2.865 6.165 3.025 ;
      RECT 6.005 2.45 6.165 3.025 ;
      RECT 6.085 1.46 6.255 2.655 ;
      RECT 3.89 2.045 5.05 2.305 ;
      RECT 4.76 0.91 4.935 2.305 ;
      RECT 6.085 1.46 6.56 1.76 ;
      RECT 4.67 0.91 4.935 1.17 ;
      RECT 5.245 2.255 5.56 2.515 ;
      RECT 5.245 0.475 5.405 2.515 ;
      RECT 2.4 1.25 2.645 1.545 ;
      RECT 2.4 1.25 2.9 1.42 ;
      RECT 2.74 0.45 2.9 1.42 ;
      RECT 5.15 0.475 5.435 1.31 ;
      RECT 3.65 1.105 4.49 1.265 ;
      RECT 4.33 0.475 4.49 1.265 ;
      RECT 3.65 0.45 3.81 1.265 ;
      RECT 4.33 0.475 5.435 0.645 ;
      RECT 2.74 0.45 3.81 0.61 ;
      RECT 3.39 1.5 3.65 2.935 ;
      RECT 3.305 1.315 3.47 1.935 ;
      RECT 3.305 1.5 4.575 1.72 ;
      RECT 3.195 0.79 3.37 1.47 ;
      RECT 3.08 0.79 3.37 0.99 ;
      RECT 1.25 2.56 1.51 3.14 ;
      RECT 2.88 2.175 3.14 2.935 ;
      RECT 1.25 2.595 3.14 2.76 ;
      RECT 1.25 2.56 1.87 2.76 ;
      RECT 1.71 1.52 1.87 2.76 ;
      RECT 0.97 1.52 1.87 1.68 ;
      RECT 0.97 0.755 1.14 1.68 ;
      RECT 0.74 0.755 1.14 1.18 ;
      RECT 0.74 0.755 2.56 0.92 ;
      RECT 2.34 0.655 2.56 0.92 ;
      RECT 2.335 1.765 2.635 2.37 ;
      RECT 2.05 1.765 3.125 1.935 ;
      RECT 2.835 1.64 3.125 1.935 ;
      RECT 2.05 1.1 2.22 1.935 ;
      RECT 1.82 1.1 2.22 1.34 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_slgcp_1

MACRO sg13g2_tiehi
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_tiehi 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.135 3.095 0.395 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.76 -0.22 1.02 0.76 ;
    END
  END VSS
  PIN L_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3927 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 2.165 1.585 2.91 ;
    END
  END L_HI
  OBS
    LAYER Metal1 ;
      RECT 0.135 2.19 0.395 2.45 ;
      RECT 0.195 1.815 0.395 2.45 ;
      RECT 0.195 1.815 1.12 2.03 ;
      RECT 0.87 1.355 1.12 2.03 ;
      RECT 1.3 0.985 1.575 1.955 ;
      RECT 0.135 0.995 0.395 1.635 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_tiehi

MACRO sg13g2_tielo
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_tielo 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.455 3.165 0.78 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.465 -0.22 0.815 0.605 ;
    END
  END VSS
  PIN L_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.295 0.485 1.585 1.23 ;
        RECT 1.095 0.485 1.585 0.775 ;
    END
  END L_LO
  OBS
    LAYER Metal1 ;
      RECT 0.875 1.03 1.115 2.06 ;
      RECT 0.315 1.03 1.115 1.29 ;
      RECT 1.305 1.46 1.58 2.875 ;
      RECT 0.315 2.11 0.575 2.76 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_tielo

MACRO sg13g2_xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_xnor2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7332 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.67 2.08 3.57 2.24 ;
        RECT 3.41 0.61 3.57 2.24 ;
        RECT 3.315 0.61 3.57 1.21 ;
        RECT 2.67 2.08 3 3.16 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4342 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.76 1.525 2.075 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4342 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.32 1.605 2.635 1.865 ;
        RECT 1.42 2.08 2.48 2.24 ;
        RECT 2.32 1.605 2.48 2.24 ;
        RECT 1.42 1.525 1.58 2.24 ;
        RECT 1.24 1.525 1.58 1.9 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.18 2.56 3.44 4 ;
        RECT 1.725 2.56 1.985 4 ;
        RECT 0.32 2.365 0.58 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.265 -0.22 2.525 0.65 ;
        RECT 0.32 -0.22 0.585 1.42 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.02 2.365 1.28 2.965 ;
      RECT 0.8 2.365 1.28 2.565 ;
      RECT 0.8 0.835 0.96 2.565 ;
      RECT 2.93 1.555 3.23 1.815 ;
      RECT 2.93 1.18 3.1 1.815 ;
      RECT 1.21 1.18 3.1 1.34 ;
      RECT 1.21 0.835 1.47 1.34 ;
      RECT 0.8 0.835 1.47 0.995 ;
      RECT 1.725 0.83 3.065 1 ;
      RECT 2.77 0.79 3.065 1 ;
      RECT 1.725 0.8 2.025 1 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_xnor2_1

MACRO sg13g2_xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_xor2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4433 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.53 1.55 2.89 1.83 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4433 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 1.55 0.82 1.83 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7064 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.45 2.155 3.71 3.16 ;
        RECT 3.53 1.115 3.71 3.16 ;
        RECT 2.835 1.115 3.71 1.315 ;
        RECT 2.835 0.67 3.1 1.315 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.43 2.9 2.69 4 ;
        RECT 0.435 2.22 0.695 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.37 -0.22 3.63 0.935 ;
        RECT 1.9 -0.22 2.16 1.27 ;
        RECT 0.285 -0.22 0.82 1.12 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.32 2.17 1.58 3.16 ;
      RECT 1.03 2.17 3.27 2.34 ;
      RECT 3.11 1.57 3.27 2.34 ;
      RECT 1.03 0.86 1.2 2.34 ;
      RECT 3.11 1.57 3.35 1.83 ;
      RECT 1.03 0.86 1.365 1.12 ;
      RECT 2.94 2.52 3.2 3.16 ;
      RECT 1.92 2.52 2.18 3.16 ;
      RECT 1.92 2.52 3.2 2.68 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_xor2_1

END LIBRARY
